module sha2_top (
    input clk,
    input rst,
    input [31:0] din,
    output [31:0] dout,
    output src_read,
    input src_ready,
    input dst_ready,
    output dst_write
);


  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire [31:0] _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire [31:0] _023_;
  wire [31:0] _024_;
  wire [31:0] _025_;
  wire [31:0] _026_;
  wire [31:0] _027_;
  wire [31:0] _028_;
  wire [31:0] _029_;
  wire [31:0] _030_;
  wire [31:0] _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire [31:0] _035_;
  wire [31:0] _036_;
  wire [31:0] _037_;
  wire [31:0] _038_;
  wire [31:0] _039_;
  wire [31:0] _040_;
  wire [31:0] _041_;
  wire [31:0] _042_;
  wire [31:0] _043_;
  wire [31:0] _044_;
  wire [31:0] _045_;
  wire [31:0] _046_;
  wire [31:0] _047_;
  wire [31:0] _048_;
  wire [31:0] _049_;
  wire [31:0] _050_;
  wire [31:0] _051_;
  wire [31:0] _052_;
  wire [31:0] _053_;
  wire [31:0] _054_;
  wire _055_;
  wire [31:0] _056_;
  wire [31:0] _057_;
  wire [31:0] _058_;
  wire [31:0] _059_;
  wire [31:0] _060_;
  wire [31:0] _061_;
  wire [31:0] _062_;
  wire [31:0] _063_;
  wire [31:0] _064_;
  wire [31:0] _065_;
  wire [31:0] _066_;
  wire [31:0] _067_;
  wire [31:0] _068_;
  wire [31:0] _069_;
  wire [31:0] _070_;
  wire [31:0] _071_;
  wire [5:0] _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire [3:0] _077_;
  wire [31:0] _078_;
  wire [21:0] _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  reg _093_;
  wire _094_;
  wire _095_;
  reg _096_;
  wire _097_;
  wire _098_;
  reg _099_;
  wire [5:0] _100_;
  wire [2047:0] _101_;
  wire [31:0] _102_;
  wire [31:0] _103_;
  wire [31:0] _104_;
  wire [31:0] _105_;
  wire [31:0] _106_;
  wire [31:0] _107_;
  wire [31:0] _108_;
  wire [31:0] _109_;
  wire [31:0] _110_;
  wire [31:0] _111_;
  reg [31:0] _112_;
  wire [31:0] _113_;
  reg [31:0] _114_;
  wire [31:0] _115_;
  reg [31:0] _116_;
  wire [31:0] _117_;
  reg [31:0] _118_;
  wire [31:0] _119_;
  reg [31:0] _120_;
  wire [31:0] _121_;
  reg [31:0] _122_;
  wire [31:0] _123_;
  reg [31:0] _124_;
  wire [31:0] _125_;
  reg [31:0] _126_;
  wire [31:0] _127_;
  reg [31:0] _128_;
  wire [31:0] _129_;
  reg [31:0] _130_;
  wire [31:0] _131_;
  reg [31:0] _132_;
  wire [31:0] _133_;
  reg [31:0] _134_;
  wire [31:0] _135_;
  reg [31:0] _136_;
  wire [31:0] _137_;
  reg [31:0] _138_;
  wire [31:0] _139_;
  reg [31:0] _140_;
  wire [31:0] _141_;
  reg [31:0] _142_;
  wire [31:0] _143_;
  wire [31:0] _144_;
  wire [31:0] _145_;
  wire [31:0] _146_;
  wire [31:0] _147_;
  wire [31:0] _148_;
  reg [31:0] _149_;
  wire [31:0] _150_;
  wire [31:0] _151_;
  reg [31:0] _152_;
  wire [21:0] _153_;
  wire [21:0] _154_;
  wire _155_;
  wire [21:0] _156_;
  wire [21:0] _157_;
  reg [21:0] _158_;
  wire [31:0] _159_;
  wire [31:0] _160_;
  reg [31:0] _161_;
  wire [31:0] _162_;
  wire [31:0] _163_;
  reg [31:0] _164_;
  wire [31:0] _165_;
  wire [31:0] _166_;
  reg [31:0] _167_;
  wire [31:0] _168_;
  wire [31:0] _169_;
  reg [31:0] _170_;
  wire [31:0] _171_;
  wire [31:0] _172_;
  reg [31:0] _173_;
  wire [31:0] _174_;
  wire [31:0] _175_;
  reg [31:0] _176_;
  wire [31:0] _177_;
  wire [31:0] _178_;
  reg [31:0] _179_;
  wire [31:0] _180_;
  wire [31:0] _181_;
  reg [31:0] _182_;
  wire [31:0] _183_;
  wire [31:0] _184_;
  reg [31:0] _185_;
  wire _186_;
  wire [3:0] _187_;
  wire [3:0] _188_;
  wire [3:0] _189_;
  reg [3:0] _190_;
  wire _191_;
  wire [5:0] _192_;
  wire [5:0] _193_;
  wire [5:0] _194_;
  reg [5:0] _195_;
  wire [31:0] _196_;
  wire [31:0] _197_;
  wire [31:0] _198_;
  wire [31:0] _199_;
  wire [31:0] _200_;
  wire [31:0] _201_;
  wire [31:0] _202_;
  wire [31:0] _203_;
  wire [31:0] _204_;
  wire [31:0] _205_;
  wire [31:0] _206_;
  wire [31:0] _207_;
  wire [31:0] _208_;
  wire [31:0] _209_;
  wire [31:0] _210_;
  wire [31:0] _211_;
  wire [31:0] _212_;
  wire [31:0] _213_;
  wire [31:0] _214_;
  wire [31:0] _215_;
  wire [31:0] _216_;
  wire [31:0] _217_;
  wire [31:0] _218_;
  wire [31:0] _219_;
  wire [31:0] _220_;
  wire [31:0] _221_;
  wire [31:0] _222_;
  wire [31:0] _223_;
  wire [31:0] _224_;
  reg [31:0] _225_;
  wire [31:0] _226_;
  wire [31:0] _227_;
  reg [31:0] _228_;
  wire [31:0] _229_;
  wire [31:0] _230_;
  reg [31:0] _231_;
  wire [31:0] _232_;
  wire [31:0] _233_;
  reg [31:0] _234_;
  wire [31:0] _235_;
  wire [31:0] _236_;
  reg [31:0] _237_;
  wire [31:0] _238_;
  wire [31:0] _239_;
  reg [31:0] _240_;
  wire [31:0] _241_;
  wire [31:0] _242_;
  reg [31:0] _243_;
  wire [31:0] _244_;
  wire [31:0] _245_;
  reg [31:0] _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire _350_;
  wire _351_;
  wire _352_;
  wire _353_;
  wire _354_;
  wire _355_;
  wire _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire _360_;
  wire _361_;
  wire _362_;
  wire _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire _367_;
  wire _368_;
  wire _369_;
  wire _370_;
  wire _371_;
  wire _372_;
  wire _373_;
  wire _374_;
  wire _375_;
  wire _376_;
  wire _377_;
  wire _378_;
  wire _379_;
  wire _380_;
  wire _381_;
  wire _382_;
  wire _383_;
  wire _384_;
  wire _385_;
  wire _386_;
  wire [4:0] _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire _391_;
  reg [4:0] _392_;
  wire _393_;
  wire [4:0] _394_;
  wire _395_;
  wire _396_;
  wire _397_;
  wire [4:0] _398_;
  wire _399_;
  wire [4:0] _400_;
  wire _401_;
  wire [4:0] _402_;
  wire _403_;
  wire [4:0] _404_;
  wire _405_;
  wire _406_;
  wire [4:0] _407_;
  wire _408_;
  wire [4:0] _409_;
  wire _410_;
  wire [4:0] _411_;
  wire _412_;
  wire [4:0] _413_;
  wire _414_;
  wire _415_;
  wire _416_;
  wire _417_;
  wire _418_;
  wire [4:0] _419_;
  wire _420_;
  wire _421_;
  wire _422_;
  wire _423_;
  wire [4:0] _424_;
  wire [4:0] _425_;
  wire [4:0] _426_;
  wire _427_;
  wire [4:0] _428_;
  wire _429_;
  wire _430_;
  wire _431_;
  wire [4:0] _432_;
  wire _433_;
  wire _434_;
  wire _435_;
  wire [4:0] _436_;
  wire _437_;
  wire _438_;
  wire _439_;
  wire _440_;
  wire _441_;
  wire _442_;
  wire _443_;
  wire _444_;
  wire _445_;
  wire _446_;
  wire _447_;
  wire _448_;
  wire _449_;
  wire _450_;
  wire _451_;
  wire _452_;
  wire _453_;
  wire _454_;
  wire _455_;
  wire _456_;
  wire _457_;
  wire _458_;
  wire _459_;
  wire _460_;
  wire _461_;
  wire _462_;
  wire _463_;
  wire _464_;
  wire _465_;
  wire _466_;
  wire _467_;
  
  wire ctr_ena_reg;
  wire ctrl_rst_reg;
  wire \dp256_gen.datapath.bf.clk ;
  wire \dp256_gen.datapath.bf.en ;
  wire [31:0] \dp256_gen.datapath.bf.exam_block ;
  wire \dp256_gen.datapath.bf.last_block_in ;
  wire \dp256_gen.datapath.bf.last_block_out ;
  wire \dp256_gen.datapath.bf.o8 ;
  wire \dp256_gen.datapath.bf.o8_in ;
  wire [3:0] \dp256_gen.datapath.bf.out_ctr ;
  wire \dp256_gen.datapath.bf.r0.clk ;
  wire \dp256_gen.datapath.bf.r0.d ;
  wire \dp256_gen.datapath.bf.r0.ena ;
  wire \dp256_gen.datapath.bf.r0.q ;
  wire \dp256_gen.datapath.bf.r0.r ;
  wire \dp256_gen.datapath.bf.r0.rst ;
  wire \dp256_gen.datapath.bf.r0:979 ;
  wire \dp256_gen.datapath.bf.r1.clk ;
  wire \dp256_gen.datapath.bf.r1.d ;
  wire \dp256_gen.datapath.bf.r1.ena ;
  wire \dp256_gen.datapath.bf.r1.q ;
  wire \dp256_gen.datapath.bf.r1.r ;
  wire \dp256_gen.datapath.bf.r1.rst ;
  wire \dp256_gen.datapath.bf.r1:982 ;
  wire \dp256_gen.datapath.bf.r4.clk ;
  wire \dp256_gen.datapath.bf.r4.d ;
  wire \dp256_gen.datapath.bf.r4.ena ;
  wire \dp256_gen.datapath.bf.r4.q ;
  wire \dp256_gen.datapath.bf.r4.r ;
  wire \dp256_gen.datapath.bf.r4.rst ;
  wire \dp256_gen.datapath.bf.r4:985 ;
  wire [5:0] \dp256_gen.datapath.bf.rd_num ;
  wire \dp256_gen.datapath.bf.rst ;
  wire \dp256_gen.datapath.bf.rst_flags ;
  wire \dp256_gen.datapath.bf.wr_len ;
  wire \dp256_gen.datapath.bf.z16 ;
  wire \dp256_gen.datapath.bf.z16_in ;
  wire \dp256_gen.datapath.bf.z16_out ;
  wire \dp256_gen.datapath.bf.zlast ;
  wire \dp256_gen.datapath.bf.zlast_in ;
  wire \dp256_gen.datapath.bf.zlast_out ;
  wire [21:0] \dp256_gen.datapath.chunk_ctr ;
  wire \dp256_gen.datapath.clk ;
  wire [5:0] \dp256_gen.datapath.const.address ;
  wire [31:0] \dp256_gen.datapath.const.output ;
  wire \dp256_gen.datapath.ctr_ena ;
  wire [31:0] \dp256_gen.datapath.data ;
  wire [31:0] \dp256_gen.datapath.dataout ;
  wire [31:0] \dp256_gen.datapath.dc.a32.d0.o ;
  wire [2:0] \dp256_gen.datapath.dc.a32.d0.tmp ;
  wire [31:0] \dp256_gen.datapath.dc.a32.d0.x ;
  wire [31:0] \dp256_gen.datapath.dc.a32.d1.o ;
  wire [9:0] \dp256_gen.datapath.dc.a32.d1.tmp ;
  wire [31:0] \dp256_gen.datapath.dc.a32.d1.x ;
  wire \dp256_gen.datapath.dc.clk ;
  wire [31:0] \dp256_gen.datapath.dc.d_one_wire ;
  wire [31:0] \dp256_gen.datapath.dc.d_zero_wire ;
  wire [31:0] \dp256_gen.datapath.dc.data ;
  wire [31:0] \dp256_gen.datapath.dc.first_stage ;
  wire \dp256_gen.datapath.dc.reg01.clk ;
  wire \dp256_gen.datapath.dc.reg01.en ;
  wire [31:0] \dp256_gen.datapath.dc.reg01.input ;
  wire [31:0] \dp256_gen.datapath.dc.reg01.output ;
  wire \dp256_gen.datapath.dc.reg01.rst ;
  wire \dp256_gen.datapath.dc.reg02.clk ;
  wire \dp256_gen.datapath.dc.reg02.en ;
  wire [31:0] \dp256_gen.datapath.dc.reg02.input ;
  wire [31:0] \dp256_gen.datapath.dc.reg02.output ;
  wire \dp256_gen.datapath.dc.reg02.rst ;
  wire [31:0] \dp256_gen.datapath.dc.second_stage ;
  wire \dp256_gen.datapath.dc.sel ;
  wire [31:0] \dp256_gen.datapath.dc.to_second_stage ;
  wire [31:0] \dp256_gen.datapath.dc.to_third_stage ;
  wire [31:0] \dp256_gen.datapath.dc.w ;
  wire [543:0] \dp256_gen.datapath.dc.wires ;
  wire \dp256_gen.datapath.dc.wr_data ;
  wire [31:0] \dp256_gen.datapath.dc.wwires ;
  wire \dp256_gen.datapath.decounter_gen.clk ;
  wire \dp256_gen.datapath.decounter_gen.ctrl ;
  wire \dp256_gen.datapath.decounter_gen.en ;
  wire [21:0] \dp256_gen.datapath.decounter_gen.input ;
  wire \dp256_gen.datapath.decounter_gen.load ;
  wire [21:0] \dp256_gen.datapath.decounter_gen.output ;
  wire [21:0] \dp256_gen.datapath.decounter_gen.reg_in ;
  wire [21:0] \dp256_gen.datapath.decounter_gen.reg_out ;
  wire \dp256_gen.datapath.decounter_gen.rst ;
  wire [21:0] \dp256_gen.datapath.decounter_gen:603 ;
  wire \dp256_gen.datapath.dst_write ;
  wire \dp256_gen.datapath.ena_reg ;
  wire [255:0] \dp256_gen.datapath.from_final_add ;
  wire [255:0] \dp256_gen.datapath.from_mux ;
  wire [255:0] \dp256_gen.datapath.from_round ;
  wire [1:0] \dp256_gen.datapath.gh ;
  wire [31:0] \dp256_gen.datapath.h_exception ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.clk ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.en ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.input ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.output ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.rst ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:1.rr:561 ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.clk ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.en ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.input ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.output ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.rst ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:2.rr:565 ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.clk ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.en ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.input ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.output ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.rst ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:3.rr:569 ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.clk ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.en ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.input ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.output ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.rst ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:4.rr:573 ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.clk ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.en ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.input ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.output ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.rst ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:5.rr:577 ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.clk ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.en ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.input ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.output ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.rst ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:6.rr:581 ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.clk ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.en ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.input ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.output ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.rst ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:7.rr:585 ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.clk ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.en ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.input ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.output ;
  wire \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.rst ;
  wire [31:0] \dp256_gen.datapath.hs256_gen.rr_gen:8.rr:589 ;
  wire \dp256_gen.datapath.kw_wr ;
  wire \dp256_gen.datapath.kwh_reg.clk ;
  wire \dp256_gen.datapath.kwh_reg.en ;
  wire [31:0] \dp256_gen.datapath.kwh_reg.input ;
  wire [31:0] \dp256_gen.datapath.kwh_reg.output ;
  wire \dp256_gen.datapath.kwh_reg.rst ;
  wire [31:0] \dp256_gen.datapath.kwh_reg:469 ;
  wire [31:0] \dp256_gen.datapath.kwhreg ;
  wire [31:0] \dp256_gen.datapath.kwhwire ;
  wire [31:0] \dp256_gen.datapath.kwire ;
  wire \dp256_gen.datapath.last_block ;
  wire \dp256_gen.datapath.last_block_out ;
  wire \dp256_gen.datapath.msg_done ;
  wire \dp256_gen.datapath.o8 ;
  wire \dp256_gen.datapath.o_ctr.clk ;
  wire [3:0] \dp256_gen.datapath.o_ctr.ctr ;
  wire \dp256_gen.datapath.o_ctr.ena ;
  wire [3:0] \dp256_gen.datapath.o_ctr.reg ;
  wire \dp256_gen.datapath.o_ctr.reset ;
  wire [3:0] \dp256_gen.datapath.out_ctr ;
  wire \dp256_gen.datapath.rd_ctr.clk ;
  wire [5:0] \dp256_gen.datapath.rd_ctr.ctr ;
  wire \dp256_gen.datapath.rd_ctr.ena ;
  wire [5:0] \dp256_gen.datapath.rd_ctr.reg ;
  wire \dp256_gen.datapath.rd_ctr.reset ;
  wire [5:0] \dp256_gen.datapath.rd_num ;
  wire [255:0] \dp256_gen.datapath.result ;
  wire [31:0] \dp256_gen.datapath.round.a32.s0.o ;
  wire [21:0] \dp256_gen.datapath.round.a32.s0.tmp ;
  wire [31:0] \dp256_gen.datapath.round.a32.s0.x ;
  wire [31:0] \dp256_gen.datapath.round.a32.s1.o ;
  wire [24:0] \dp256_gen.datapath.round.a32.s1.tmp ;
  wire [31:0] \dp256_gen.datapath.round.a32.s1.x ;
  wire [31:0] \dp256_gen.datapath.round.ain ;
  wire [31:0] \dp256_gen.datapath.round.aout ;
  wire [31:0] \dp256_gen.datapath.round.bin ;
  wire [31:0] \dp256_gen.datapath.round.bout ;
  wire [31:0] \dp256_gen.datapath.round.c1.o ;
  wire [31:0] \dp256_gen.datapath.round.c1.x ;
  wire [31:0] \dp256_gen.datapath.round.c1.y ;
  wire [31:0] \dp256_gen.datapath.round.c1.z ;
  wire [31:0] \dp256_gen.datapath.round.cf0_reg ;
  wire [31:0] \dp256_gen.datapath.round.cf1_reg ;
  wire [31:0] \dp256_gen.datapath.round.ch_reg ;
  wire [31:0] \dp256_gen.datapath.round.cin ;
  wire [31:0] \dp256_gen.datapath.round.cout ;
  wire [31:0] \dp256_gen.datapath.round.din ;
  wire [31:0] \dp256_gen.datapath.round.dout ;
  wire [31:0] \dp256_gen.datapath.round.ein ;
  wire [31:0] \dp256_gen.datapath.round.eout ;
  wire [31:0] \dp256_gen.datapath.round.fin ;
  wire [31:0] \dp256_gen.datapath.round.fout ;
  wire [31:0] \dp256_gen.datapath.round.g_or_h ;
  wire [31:0] \dp256_gen.datapath.round.gin ;
  wire [31:0] \dp256_gen.datapath.round.gout ;
  wire [31:0] \dp256_gen.datapath.round.hin ;
  wire [31:0] \dp256_gen.datapath.round.hout ;
  wire [31:0] \dp256_gen.datapath.round.kw ;
  wire [31:0] \dp256_gen.datapath.round.kwhwire ;
  wire [31:0] \dp256_gen.datapath.round.kwire ;
  wire [31:0] \dp256_gen.datapath.round.m1.o ;
  wire [31:0] \dp256_gen.datapath.round.m1.x ;
  wire [31:0] \dp256_gen.datapath.round.m1.y ;
  wire [31:0] \dp256_gen.datapath.round.m1.z ;
  wire [31:0] \dp256_gen.datapath.round.maj_reg ;
  wire \dp256_gen.datapath.round.sel_gh ;
  wire [31:0] \dp256_gen.datapath.round.wwire ;
  wire \dp256_gen.datapath.rst ;
  wire \dp256_gen.datapath.rst_flags ;
  wire \dp256_gen.datapath.sel ;
  wire \dp256_gen.datapath.sel2 ;
  wire \dp256_gen.datapath.sel_gh ;
  wire \dp256_gen.datapath.sel_gh2 ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.clk ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.en ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.input ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.output ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.rst ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:1.sr0:438 ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.clk ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.en ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.input ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.output ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.rst ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:2.sr0:442 ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.clk ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.en ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.input ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.output ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.rst ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:3.sr0:446 ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.clk ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.en ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.input ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.output ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.rst ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:4.sr0:450 ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.clk ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.en ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.input ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.output ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.rst ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:5.sr0:454 ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.clk ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.en ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.input ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.output ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.rst ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:6.sr0:458 ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.clk ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.en ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.input ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.output ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.rst ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:7.sr0:462 ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.clk ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.en ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.input ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.output ;
  wire \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.rst ;
  wire [31:0] \dp256_gen.datapath.st256_gen.sr_gen:8.sr0:466 ;
  wire [255:0] \dp256_gen.datapath.to_result ;
  wire [255:0] \dp256_gen.datapath.to_round ;
  wire \dp256_gen.datapath.wr_chctr ;
  wire \dp256_gen.datapath.wr_data ;
  wire \dp256_gen.datapath.wr_len ;
  wire \dp256_gen.datapath.wr_result ;
  wire \dp256_gen.datapath.wr_state ;
  wire [31:0] \dp256_gen.datapath.wwire ;
  wire \dp256_gen.datapath.z16 ;
  wire \dp256_gen.datapath.z16_reg ;
  wire \dp256_gen.datapath.zlast ;
  wire dst_write_reg;
  wire kr_wr_wire;
  wire lb_reg;
  wire msg_done_reg;
  wire o8_reg;
  wire \rsc0.clk ;
  wire \rsc0.ctr_ena ;
  wire \rsc0.ctrl_rst ;
  wire [4:0] \rsc0.current_state ;
  wire \rsc0.dst_ready ;
  wire \rsc0.dst_write ;
  wire \rsc0.kw_wr ;
  wire \rsc0.last_block ;
  wire \rsc0.msg_done ;
  wire [4:0] \rsc0.next_state ;
  wire \rsc0.o8 ;
  wire \rsc0.rst ;
  wire \rsc0.rst_flags ;
  wire \rsc0.sel ;
  wire \rsc0.sel2 ;
  wire \rsc0.sel_gh ;
  wire \rsc0.sel_gh2 ;
  wire \rsc0.src_read ;
  wire \rsc0.src_read_sig ;
  wire \rsc0.src_ready ;
  wire \rsc0.wr_chctr ;
  wire \rsc0.wr_data ;
  wire \rsc0.wr_len ;
  wire \rsc0.wr_result ;
  wire \rsc0.wr_state ;
  wire \rsc0.z16 ;
  wire \rsc0.zlast ;
  wire rst_flags_reg;
  wire rst_reg;
  wire sel2_reg;
  wire sel_gh_reg;
  wire sel_gh_reg2;
  wire sel_reg;
  wire src_ready_reg;
  wire wr_chctr_reg;
  wire wr_data_reg;
  wire wr_len_reg;
  wire wr_result_reg;
  wire wr_state_reg;
  wire z16_reg;
  wire zlast_reg;
  reg [31:0] \dp256_gen.datapath.const.1017 [63:0];
  initial begin
    \dp256_gen.datapath.const.1017 [0]  = 32'd3329325298;
    \dp256_gen.datapath.const.1017 [1]  = 32'd3204031479;
    \dp256_gen.datapath.const.1017 [2]  = 32'd2756734187;
    \dp256_gen.datapath.const.1017 [3]  = 32'd2428436474;
    \dp256_gen.datapath.const.1017 [4]  = 32'd2361852424;
    \dp256_gen.datapath.const.1017 [5]  = 32'd2227730452;
    \dp256_gen.datapath.const.1017 [6]  = 32'd2024104815;
    \dp256_gen.datapath.const.1017 [7]  = 32'd1955562222;
    \dp256_gen.datapath.const.1017 [8]  = 32'd1747873779;
    \dp256_gen.datapath.const.1017 [9]  = 32'd1537002063;
    \dp256_gen.datapath.const.1017 [10] = 32'd1322822218;
    \dp256_gen.datapath.const.1017 [11] = 32'd958139571;
    \dp256_gen.datapath.const.1017 [12] = 32'd883997877;
    \dp256_gen.datapath.const.1017 [13] = 32'd659060556;
    \dp256_gen.datapath.const.1017 [14] = 32'd506948616;
    \dp256_gen.datapath.const.1017 [15] = 32'd430227734;
    \dp256_gen.datapath.const.1017 [16] = 32'd275423344;
    \dp256_gen.datapath.const.1017 [17] = 32'd4094571909;
    \dp256_gen.datapath.const.1017 [18] = 32'd3600352804;
    \dp256_gen.datapath.const.1017 [19] = 32'd3516065817;
    \dp256_gen.datapath.const.1017 [20] = 32'd3345764771;
    \dp256_gen.datapath.const.1017 [21] = 32'd3259730800;
    \dp256_gen.datapath.const.1017 [22] = 32'd2820302411;
    \dp256_gen.datapath.const.1017 [23] = 32'd2730485921;
    \dp256_gen.datapath.const.1017 [24] = 32'd2456956037;
    \dp256_gen.datapath.const.1017 [25] = 32'd2177026350;
    \dp256_gen.datapath.const.1017 [26] = 32'd1986661051;
    \dp256_gen.datapath.const.1017 [27] = 32'd1695183700;
    \dp256_gen.datapath.const.1017 [28] = 32'd1396182291;
    \dp256_gen.datapath.const.1017 [29] = 32'd1294757372;
    \dp256_gen.datapath.const.1017 [30] = 32'd773529912;
    \dp256_gen.datapath.const.1017 [31] = 32'd666307205;
    \dp256_gen.datapath.const.1017 [32] = 32'd338241895;
    \dp256_gen.datapath.const.1017 [33] = 32'd113926993;
    \dp256_gen.datapath.const.1017 [34] = 32'd3584528711;
    \dp256_gen.datapath.const.1017 [35] = 32'd3336571891;
    \dp256_gen.datapath.const.1017 [36] = 32'd3210313671;
    \dp256_gen.datapath.const.1017 [37] = 32'd2952996808;
    \dp256_gen.datapath.const.1017 [38] = 32'd2821834349;
    \dp256_gen.datapath.const.1017 [39] = 32'd2554220882;
    \dp256_gen.datapath.const.1017 [40] = 32'd1996064986;
    \dp256_gen.datapath.const.1017 [41] = 32'd1555081692;
    \dp256_gen.datapath.const.1017 [42] = 32'd1249150122;
    \dp256_gen.datapath.const.1017 [43] = 32'd770255983;
    \dp256_gen.datapath.const.1017 [44] = 32'd604807628;
    \dp256_gen.datapath.const.1017 [45] = 32'd264347078;
    \dp256_gen.datapath.const.1017 [46] = 32'd4022224774;
    \dp256_gen.datapath.const.1017 [47] = 32'd3835390401;
    \dp256_gen.datapath.const.1017 [48] = 32'd3248222580;
    \dp256_gen.datapath.const.1017 [49] = 32'd2614888103;
    \dp256_gen.datapath.const.1017 [50] = 32'd2162078206;
    \dp256_gen.datapath.const.1017 [51] = 32'd1925078388;
    \dp256_gen.datapath.const.1017 [52] = 32'd1426881987;
    \dp256_gen.datapath.const.1017 [53] = 32'd607225278;
    \dp256_gen.datapath.const.1017 [54] = 32'd310598401;
    \dp256_gen.datapath.const.1017 [55] = 32'd3624381080;
    \dp256_gen.datapath.const.1017 [56] = 32'd2870763221;
    \dp256_gen.datapath.const.1017 [57] = 32'd2453635748;
    \dp256_gen.datapath.const.1017 [58] = 32'd1508970993;
    \dp256_gen.datapath.const.1017 [59] = 32'd961987163;
    \dp256_gen.datapath.const.1017 [60] = 32'd3921009573;
    \dp256_gen.datapath.const.1017 [61] = 32'd3049323471;
    \dp256_gen.datapath.const.1017 [62] = 32'd1899447441;
    \dp256_gen.datapath.const.1017 [63] = 32'd1116352408;
  end
  assign _102_ = \dp256_gen.datapath.const.1017 [_100_];
  assign _000_ = ~src_ready;
  assign _011_ = ctrl_rst_reg | rst;
  assign _032_ = !\dp256_gen.datapath.gh ;
  assign _033_ = \dp256_gen.datapath.gh == 2'h1;
  assign _034_ = \dp256_gen.datapath.gh == 2'h2;
  function [31:0] \dp256_gen.datapath.484 ;
    input [31:0] a;
    input [95:0] b;
    input [2:0] s;
    casez (s)  // synopsys parallel_case
      3'b??1:  \dp256_gen.datapath.484 = b[31:0];
      3'b?1?:  \dp256_gen.datapath.484 = b[63:32];
      3'b1??:  \dp256_gen.datapath.484 = b[95:64];
      default: \dp256_gen.datapath.484 = a;
    endcase
  endfunction
  assign _035_ = \dp256_gen.datapath.484 (
      \dp256_gen.datapath.result [63:32],
      {
        \dp256_gen.datapath.to_round [31:0], \dp256_gen.datapath.to_round [63:32], \dp256_gen.datapath.to_round [63:32]
      },
      {
        _034_, _033_, _032_
      }
  );
  assign _045_ = \dp256_gen.datapath.to_round [255:224] + \dp256_gen.datapath.result [159:128];
  assign _046_ = \dp256_gen.datapath.to_round [127:96] + \dp256_gen.datapath.result [31:0];
  assign _047_ = \dp256_gen.datapath.sel  ? \dp256_gen.datapath.from_final_add [255:224] : \dp256_gen.datapath.from_round [255:224];
  assign _048_ = \dp256_gen.datapath.sel  ? \dp256_gen.datapath.from_final_add [223:192] : \dp256_gen.datapath.from_round [223:192];
  assign _049_ = \dp256_gen.datapath.sel  ? \dp256_gen.datapath.from_final_add [191:160] : \dp256_gen.datapath.from_round [191:160];
  assign _050_ = \dp256_gen.datapath.sel  ? \dp256_gen.datapath.from_final_add [159:128] : \dp256_gen.datapath.from_round [159:128];
  assign _051_ = \dp256_gen.datapath.sel  ? \dp256_gen.datapath.from_final_add [127:96] : \dp256_gen.datapath.from_round [127:96];
  assign _052_ = \dp256_gen.datapath.sel  ? \dp256_gen.datapath.from_final_add [95:64] : \dp256_gen.datapath.from_round [95:64];
  assign _053_ = \dp256_gen.datapath.sel  ? \dp256_gen.datapath.from_final_add [63:32] : \dp256_gen.datapath.from_round [63:32];
  assign _054_ = \dp256_gen.datapath.sel  ? \dp256_gen.datapath.from_final_add [31:0] : \dp256_gen.datapath.from_round [31:0];
  assign _055_ = \dp256_gen.datapath.wr_result | \dp256_gen.datapath.dst_write ;
  assign _056_ = \dp256_gen.datapath.wr_result  ? \dp256_gen.datapath.from_final_add [255:224] : \dp256_gen.datapath.result [223:192];
  assign _057_ = \dp256_gen.datapath.wr_result  ? \dp256_gen.datapath.from_final_add [223:192] : \dp256_gen.datapath.result [191:160];
  assign _058_ = \dp256_gen.datapath.wr_result  ? \dp256_gen.datapath.from_final_add [191:160] : \dp256_gen.datapath.result [159:128];
  assign _059_ = \dp256_gen.datapath.wr_result  ? \dp256_gen.datapath.from_final_add [159:128] : \dp256_gen.datapath.result [127:96];
  assign _060_ = \dp256_gen.datapath.wr_result  ? \dp256_gen.datapath.from_final_add [127:96] : \dp256_gen.datapath.result [95:64];
  assign _061_ = \dp256_gen.datapath.wr_result  ? \dp256_gen.datapath.from_final_add [95:64] : \dp256_gen.datapath.result [63:32];
  assign _062_ = \dp256_gen.datapath.wr_result  ? \dp256_gen.datapath.from_final_add [63:32] : \dp256_gen.datapath.result [31:0];
  assign _080_ = !\dp256_gen.datapath.chunk_ctr ;
  assign _081_ = _080_ ? 1'h1 : 1'h0;
  assign _082_ = \dp256_gen.datapath.bf.rd_num == 6'h0b;
  assign _083_ = _082_ ? 1'h1 : 1'h0;
  assign _084_ = \dp256_gen.datapath.bf.rd_num == 6'h3b;
  assign _085_ = _084_ ? 1'h1 : 1'h0;
  assign _086_ = \dp256_gen.datapath.bf.out_ctr == 4'h7;
  assign _087_ = _086_ ? 1'h1 : 1'h0;
  assign _091_ = \dp256_gen.datapath.bf.r0.ena ? \dp256_gen.datapath.bf.r0.d : \dp256_gen.datapath.bf.r0.r ;
  assign _092_ = \dp256_gen.datapath.bf.r0.rst ? 1'h0 : _091_;
  always @(posedge \dp256_gen.datapath.bf.r0.clk ) _093_ <= _092_;
  assign _094_ = \dp256_gen.datapath.bf.r1.ena ? \dp256_gen.datapath.bf.r1.d : \dp256_gen.datapath.bf.r1.r ;
  assign _095_ = \dp256_gen.datapath.bf.r1.rst ? 1'h0 : _094_;
  always @(posedge \dp256_gen.datapath.bf.r1.clk ) _096_ <= _095_;
  assign _097_ = \dp256_gen.datapath.bf.r4.ena ? \dp256_gen.datapath.bf.r4.d : \dp256_gen.datapath.bf.r4.r ;
  assign _098_ = \dp256_gen.datapath.bf.r4.rst ? 1'h0 : _097_;
  always @(posedge \dp256_gen.datapath.bf.r4.clk ) _099_ <= _098_;
  assign _100_ = 6'h3f - \dp256_gen.datapath.const.address ;
  assign _103_ = \dp256_gen.datapath.dc.sel ? \dp256_gen.datapath.dc.wwires : \dp256_gen.datapath.dc.data ;
  assign _106_ = \dp256_gen.datapath.dc.d_zero_wire + \dp256_gen.datapath.dc.wires [95:64];
  assign _108_ = \dp256_gen.datapath.dc.to_second_stage + \dp256_gen.datapath.dc.wires [351:320];
  assign _110_ = \dp256_gen.datapath.dc.to_third_stage + \dp256_gen.datapath.dc.d_one_wire ;
  assign _111_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [63:32] : \dp256_gen.datapath.dc.wires [31:0];
  always @(posedge \dp256_gen.datapath.dc.clk ) _112_ <= _111_;
  assign _113_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [95:64] : \dp256_gen.datapath.dc.wires [63:32];
  always @(posedge \dp256_gen.datapath.dc.clk ) _114_ <= _113_;
  assign _115_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [127:96] : \dp256_gen.datapath.dc.wires [95:64];
  always @(posedge \dp256_gen.datapath.dc.clk ) _116_ <= _115_;
  assign _117_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [159:128] : \dp256_gen.datapath.dc.wires [127:96];
  always @(posedge \dp256_gen.datapath.dc.clk ) _118_ <= _117_;
  assign _119_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [191:160] : \dp256_gen.datapath.dc.wires [159:128];
  always @(posedge \dp256_gen.datapath.dc.clk ) _120_ <= _119_;
  assign _121_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [223:192] : \dp256_gen.datapath.dc.wires [191:160];
  always @(posedge \dp256_gen.datapath.dc.clk ) _122_ <= _121_;
  assign _123_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [255:224] : \dp256_gen.datapath.dc.wires [223:192];
  always @(posedge \dp256_gen.datapath.dc.clk ) _124_ <= _123_;
  assign _125_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [287:256] : \dp256_gen.datapath.dc.wires [255:224];
  always @(posedge \dp256_gen.datapath.dc.clk ) _126_ <= _125_;
  assign _127_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [319:288] : \dp256_gen.datapath.dc.wires [287:256];
  always @(posedge \dp256_gen.datapath.dc.clk ) _128_ <= _127_;
  assign _129_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [351:320] : \dp256_gen.datapath.dc.wires [319:288];
  always @(posedge \dp256_gen.datapath.dc.clk ) _130_ <= _129_;
  assign _131_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [383:352] : \dp256_gen.datapath.dc.wires [351:320];
  always @(posedge \dp256_gen.datapath.dc.clk ) _132_ <= _131_;
  assign _133_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [415:384] : \dp256_gen.datapath.dc.wires [383:352];
  always @(posedge \dp256_gen.datapath.dc.clk ) _134_ <= _133_;
  assign _135_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [447:416] : \dp256_gen.datapath.dc.wires [415:384];
  always @(posedge \dp256_gen.datapath.dc.clk ) _136_ <= _135_;
  assign _137_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [479:448] : \dp256_gen.datapath.dc.wires [447:416];
  always @(posedge \dp256_gen.datapath.dc.clk ) _138_ <= _137_;
  assign _139_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [511:480] : \dp256_gen.datapath.dc.wires [479:448];
  always @(posedge \dp256_gen.datapath.dc.clk ) _140_ <= _139_;
  assign _141_ = \dp256_gen.datapath.dc.wr_data  ? \dp256_gen.datapath.dc.wires [543:512] : \dp256_gen.datapath.dc.wires [511:480];
  always @(posedge \dp256_gen.datapath.dc.clk ) _142_ <= _141_;
  assign _143_ = { \dp256_gen.datapath.dc.a32.d0.x [6:0], \dp256_gen.datapath.dc.a32.d0.x [31:7] } ^ { \dp256_gen.datapath.dc.a32.d0.x [17:0], \dp256_gen.datapath.dc.a32.d0.x [31:18] };
  assign _144_ = _143_ ^ {\dp256_gen.datapath.dc.a32.d0.tmp , \dp256_gen.datapath.dc.a32.d0.x [31:3]};
  assign _145_ = { \dp256_gen.datapath.dc.a32.d1.x [16:0], \dp256_gen.datapath.dc.a32.d1.x [31:17] } ^ { \dp256_gen.datapath.dc.a32.d1.x [18:0], \dp256_gen.datapath.dc.a32.d1.x [31:19] };
  assign _146_ = _145_ ^ {\dp256_gen.datapath.dc.a32.d1.tmp , \dp256_gen.datapath.dc.a32.d1.x [31:10]};
  assign _147_ = \dp256_gen.datapath.dc.reg01.en ? \dp256_gen.datapath.dc.reg01.input : _149_;
  assign _148_ = \dp256_gen.datapath.dc.reg01.rst ? 32'd0 : _147_;
  always @(posedge \dp256_gen.datapath.dc.reg01.clk ) _149_ <= _148_;
  assign _150_ = \dp256_gen.datapath.dc.reg02.en ? \dp256_gen.datapath.dc.reg02.input : _152_;
  assign _151_ = \dp256_gen.datapath.dc.reg02.rst ? 32'd0 : _150_;
  always @(posedge \dp256_gen.datapath.dc.reg02.clk ) _152_ <= _151_;
  assign _153_ = \dp256_gen.datapath.decounter_gen.load ? \dp256_gen.datapath.decounter_gen.input : _154_;
  assign _154_ = \dp256_gen.datapath.decounter_gen.reg_out - 22'h000001;
  assign _155_ = \dp256_gen.datapath.decounter_gen.load | \dp256_gen.datapath.decounter_gen.en ;
  assign _156_ = \dp256_gen.datapath.decounter_gen.ctrl  ? \dp256_gen.datapath.decounter_gen.reg_in  : \dp256_gen.datapath.decounter_gen.reg_out ;
  assign _157_ = \dp256_gen.datapath.decounter_gen.rst ? 22'h000000 : _156_;
  always @(posedge \dp256_gen.datapath.decounter_gen.clk ) _158_ <= _157_;
  assign _159_ = \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.en ? \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.input : _161_;
  assign _160_ = \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.rst ? 32'd1779033703 : _159_;
  always @(posedge \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.clk ) _161_ <= _160_;
  assign _162_ = \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.en ? \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.input : _164_;
  assign _163_ = \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.rst ? 32'd3144134277 : _162_;
  always @(posedge \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.clk ) _164_ <= _163_;
  assign _165_ = \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.en ? \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.input : _167_;
  assign _166_ = \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.rst ? 32'd1013904242 : _165_;
  always @(posedge \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.clk ) _167_ <= _166_;
  assign _168_ = \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.en ? \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.input : _170_;
  assign _169_ = \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.rst ? 32'd2773480762 : _168_;
  always @(posedge \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.clk ) _170_ <= _169_;
  assign _171_ = \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.en ? \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.input : _173_;
  assign _172_ = \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.rst ? 32'd1359893119 : _171_;
  always @(posedge \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.clk ) _173_ <= _172_;
  assign _174_ = \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.en ? \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.input : _176_;
  assign _175_ = \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.rst ? 32'd2600822924 : _174_;
  always @(posedge \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.clk ) _176_ <= _175_;
  assign _177_ = \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.en ? \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.input : _179_;
  assign _178_ = \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.rst ? 32'd528734635 : _177_;
  always @(posedge \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.clk ) _179_ <= _178_;
  assign _180_ = \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.en ? \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.input : _182_;
  assign _181_ = \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.rst ? 32'd1541459225 : _180_;
  always @(posedge \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.clk ) _182_ <= _181_;
  assign _183_ = \dp256_gen.datapath.kwh_reg.en ? \dp256_gen.datapath.kwh_reg.input : _185_;
  assign _184_ = \dp256_gen.datapath.kwh_reg.rst ? 32'd0 : _183_;
  always @(posedge \dp256_gen.datapath.kwh_reg.clk ) _185_ <= _184_;
  assign _187_ = \dp256_gen.datapath.o_ctr.reg + 4'h1;
  assign _188_ = _186_ ? 4'h0 : _187_;
  assign _189_ = \dp256_gen.datapath.o_ctr.ena ? _188_ : \dp256_gen.datapath.o_ctr.reg ;
  always @(posedge \dp256_gen.datapath.o_ctr.clk , posedge \dp256_gen.datapath.o_ctr.reset )
    if (\dp256_gen.datapath.o_ctr.reset ) _190_ <= 4'h0;
    else _190_ <= _189_;
  assign _186_ = \dp256_gen.datapath.o_ctr.reg == 4'h8;
  assign _191_ = \dp256_gen.datapath.rd_ctr.reg == 6'h3f;
  assign _192_ = \dp256_gen.datapath.rd_ctr.reg + 6'h01;
  assign _193_ = _191_ ? 6'h00 : _192_;
  assign _194_ = \dp256_gen.datapath.rd_ctr.ena ? _193_ : \dp256_gen.datapath.rd_ctr.reg ;
  always @(posedge \dp256_gen.datapath.rd_ctr.clk , posedge \dp256_gen.datapath.rd_ctr.reset )
    if (\dp256_gen.datapath.rd_ctr.reset ) _195_ <= 6'h00;
    else _195_ <= _194_;
  assign _200_ = \dp256_gen.datapath.round.ch_reg + \dp256_gen.datapath.round.cf1_reg ;
  assign _201_ = _200_ + \dp256_gen.datapath.round.kw ;
  assign _202_ = _201_ + \dp256_gen.datapath.round.din ;
  assign _203_ = \dp256_gen.datapath.round.kw + \dp256_gen.datapath.round.maj_reg ;
  assign _204_ = _203_ + \dp256_gen.datapath.round.cf0_reg ;
  assign _205_ = _204_ + \dp256_gen.datapath.round.ch_reg ;
  assign _206_ = _205_ + \dp256_gen.datapath.round.cf1_reg ;
  assign _207_ = \dp256_gen.datapath.round.sel_gh ? \dp256_gen.datapath.round.hin : \dp256_gen.datapath.round.gin ;
  assign _208_ = \dp256_gen.datapath.round.g_or_h + \dp256_gen.datapath.round.kwire ;
  assign _209_ = _208_ + \dp256_gen.datapath.round.wwire ;
  assign _210_ = { \dp256_gen.datapath.round.a32.s0.x [1:0], \dp256_gen.datapath.round.a32.s0.x [31:2] } ^ { \dp256_gen.datapath.round.a32.s0.x [12:0], \dp256_gen.datapath.round.a32.s0.x [31:13] };
  assign _211_ = _210_ ^ {\dp256_gen.datapath.round.a32.s0.tmp , \dp256_gen.datapath.round.a32.s0.x [31:22]};
  assign _212_ = { \dp256_gen.datapath.round.a32.s1.x [5:0], \dp256_gen.datapath.round.a32.s1.x [31:6] } ^ { \dp256_gen.datapath.round.a32.s1.x [10:0], \dp256_gen.datapath.round.a32.s1.x [31:11] };
  assign _213_ = _212_ ^ {\dp256_gen.datapath.round.a32.s1.tmp , \dp256_gen.datapath.round.a32.s1.x [31:25]};
  assign _214_ = \dp256_gen.datapath.round.c1.x & \dp256_gen.datapath.round.c1.y ;
  assign _215_ = ~\dp256_gen.datapath.round.c1.x ;
  assign _216_ = _215_ & \dp256_gen.datapath.round.c1.z ;
  assign _217_ = _214_ ^ _216_;
  assign _218_ = \dp256_gen.datapath.round.m1.x & \dp256_gen.datapath.round.m1.y ;
  assign _219_ = \dp256_gen.datapath.round.m1.x & \dp256_gen.datapath.round.m1.z ;
  assign _220_ = _218_ ^ _219_;
  assign _221_ = \dp256_gen.datapath.round.m1.y & \dp256_gen.datapath.round.m1.z ;
  assign _222_ = _220_ ^ _221_;
  assign _223_ = \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.en  ? \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.input  : _225_;
  assign _224_ = \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.rst ? 32'd1779033703 : _223_;
  always @(posedge \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.clk ) _225_ <= _224_;
  assign _226_ = \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.en  ? \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.input  : _228_;
  assign _227_ = \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.rst ? 32'd3144134277 : _226_;
  always @(posedge \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.clk ) _228_ <= _227_;
  assign _229_ = \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.en  ? \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.input  : _231_;
  assign _230_ = \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.rst ? 32'd1013904242 : _229_;
  always @(posedge \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.clk ) _231_ <= _230_;
  assign _232_ = \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.en  ? \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.input  : _234_;
  assign _233_ = \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.rst ? 32'd2773480762 : _232_;
  always @(posedge \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.clk ) _234_ <= _233_;
  assign _235_ = \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.en  ? \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.input  : _237_;
  assign _236_ = \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.rst ? 32'd1359893119 : _235_;
  always @(posedge \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.clk ) _237_ <= _236_;
  assign _238_ = \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.en  ? \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.input  : _240_;
  assign _239_ = \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.rst ? 32'd2600822924 : _238_;
  always @(posedge \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.clk ) _240_ <= _239_;
  assign _241_ = \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.en  ? \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.input  : _243_;
  assign _242_ = \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.rst ? 32'd528734635 : _241_;
  always @(posedge \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.clk ) _243_ <= _242_;
  assign _244_ = \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.en  ? \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.input  : _246_;
  assign _245_ = \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.rst ? 32'd1541459225 : _244_;
  always @(posedge \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.clk ) _246_ <= _245_;
  assign _414_ = \rsc0.current_state == 5'h09;
  assign _415_ = \rsc0.current_state == 5'h0a;
  assign _416_ = \rsc0.current_state == 5'h0b;
  assign _417_ = \rsc0.current_state == 5'h0c;
  assign _418_ = \rsc0.src_ready | \rsc0.msg_done ;
  assign _419_ = _418_ ? 5'h0e : 5'h0d;
  assign _420_ = \rsc0.current_state == 5'h0d;
  assign _421_ = \rsc0.msg_done & \rsc0.last_block ;
  assign _422_ = ~\rsc0.last_block ;
  assign _423_ = \rsc0.msg_done & _422_;
  assign _424_ = \rsc0.src_ready ? 5'h0f : 5'h0e;
  assign _425_ = _423_ ? 5'h11 : _424_;
  assign _426_ = _421_ ? 5'h10 : _425_;
  assign _427_ = \rsc0.current_state == 5'h0e;
  assign _428_ = \rsc0.src_ready ? 5'h06 : 5'h0f;
  assign _429_ = \rsc0.current_state == 5'h0f;
  assign _430_ = ~\rsc0.dst_ready ;
  assign _431_ = \rsc0.o8 & _430_;
  assign _432_ = _431_ ? 5'h12 : 5'h10;
  assign _433_ = \rsc0.current_state == 5'h10;
  assign _434_ = \rsc0.current_state == 5'h12;
  assign _435_ = \rsc0.current_state == 5'h11;
  function [4:0] \rsc0.149 ;
    input [4:0] a;
    input [94:0] b;
    input [18:0] s;
    casez (s)  // synopsys parallel_case
      19'b??????????????????1: \rsc0.149 = b[4:0];
      19'b?????????????????1?: \rsc0.149 = b[9:5];
      19'b????????????????1??: \rsc0.149 = b[14:10];
      19'b???????????????1???: \rsc0.149 = b[19:15];
      19'b??????????????1????: \rsc0.149 = b[24:20];
      19'b?????????????1?????: \rsc0.149 = b[29:25];
      19'b????????????1??????: \rsc0.149 = b[34:30];
      19'b???????????1???????: \rsc0.149 = b[39:35];
      19'b??????????1????????: \rsc0.149 = b[44:40];
      19'b?????????1?????????: \rsc0.149 = b[49:45];
      19'b????????1??????????: \rsc0.149 = b[54:50];
      19'b???????1???????????: \rsc0.149 = b[59:55];
      19'b??????1????????????: \rsc0.149 = b[64:60];
      19'b?????1?????????????: \rsc0.149 = b[69:65];
      19'b????1??????????????: \rsc0.149 = b[74:70];
      19'b???1???????????????: \rsc0.149 = b[79:75];
      19'b??1????????????????: \rsc0.149 = b[84:80];
      19'b?1?????????????????: \rsc0.149 = b[89:85];
      19'b1??????????????????: \rsc0.149 = b[94:90];
      default: \rsc0.149 = a;
    endcase
  endfunction
  assign _436_ = \rsc0.149 (
      5'hxx,
      {
        10'h021,
        _432_,
        _428_,
        _426_,
        _419_,
        15'h358b,
        _413_,
        _411_,
        _409_,
        _407_,
        _404_,
        _402_,
        _400_,
        _398_,
        _394_,
        _387_
      },
      {
        _435_,
        _434_,
        _433_,
        _429_,
        _427_,
        _420_,
        _417_,
        _416_,
        _415_,
        _414_,
        _412_,
        _410_,
        _408_,
        _405_,
        _403_,
        _401_,
        _399_,
        _395_,
        _393_
      }
  );
  assign _437_ = \rsc0.current_state == 5'h01;
  assign _438_ = \rsc0.src_ready & _437_;
  assign _439_ = _438_ ? 1'h1 : 1'h0;
  assign _440_ = \rsc0.current_state == 5'h03;
  assign _441_ = \rsc0.current_state == 5'h04;
  assign _442_ = _440_ | _441_;
  assign _443_ = \rsc0.current_state == 5'h05;
  assign _444_ = _442_ | _443_;
  assign _445_ = \rsc0.current_state == 5'h06;
  assign _446_ = _444_ | _445_;
  assign _447_ = \rsc0.current_state == 5'h07;
  assign _448_ = _446_ | _447_;
  assign _449_ = \rsc0.current_state == 5'h08;
  assign _450_ = _448_ | _449_;
  assign _451_ = \rsc0.current_state == 5'h0e;
  assign _452_ = _450_ | _451_;
  assign _453_ = \rsc0.current_state == 5'h0f;
  assign _454_ = _452_ | _453_;
  assign _455_ = \rsc0.current_state == 5'h0d;
  assign _456_ = ~\rsc0.msg_done ;
  assign _457_ = _456_ & _455_;
  assign _458_ = _454_ | _457_;
  assign _459_ = \rsc0.current_state == 5'h0e;
  assign _460_ = _458_ | _459_;
  assign _461_ = _460_ & \rsc0.src_ready ;
  assign _462_ = \rsc0.current_state == 5'h09;
  assign _463_ = _461_ | _462_;
  assign _464_ = \rsc0.current_state == 5'h0a;
  assign _465_ = _463_ | _464_;
  assign _466_ = \rsc0.current_state == 5'h0b;
  assign _467_ = _465_ | _466_;
  assign _247_ = \rsc0.current_state == 5'h0c;
  assign _248_ = _467_ | _247_;
  assign _249_ = _248_ ? 1'h1 : 1'h0;
  assign _250_ = \rsc0.current_state == 5'h0b;
  assign _251_ = \rsc0.current_state == 5'h0c;
  assign _252_ = _250_ | _251_;
  assign _253_ = \rsc0.current_state == 5'h0d;
  assign _254_ = \rsc0.src_ready | \rsc0.msg_done ;
  assign _255_ = _254_ & _253_;
  assign _256_ = _252_ | _255_;
  assign _257_ = \rsc0.current_state == 5'h0e;
  assign _258_ = \rsc0.src_ready | \rsc0.msg_done ;
  assign _259_ = _258_ & _257_;
  assign _260_ = _256_ | _259_;
  assign _261_ = _260_ ? 1'h1 : 1'h0;
  assign _262_ = \rsc0.current_state == 5'h01;
  assign _263_ = \rsc0.src_ready & _262_;
  assign _264_ = \rsc0.current_state == 5'h02;
  assign _265_ = \rsc0.last_block & _264_;
  assign _266_ = \rsc0.src_ready & _265_;
  assign _267_ = _263_ | _266_;
  assign _268_ = \rsc0.current_state == 5'h0d;
  assign _269_ = \rsc0.current_state == 5'h0e;
  assign _270_ = _268_ | _269_;
  assign _271_ = \rsc0.src_ready & _270_;
  assign _272_ = ~\rsc0.msg_done ;
  assign _273_ = _272_ & _271_;
  assign _274_ = _267_ | _273_;
  assign _275_ = \rsc0.current_state == 5'h03;
  assign _276_ = \rsc0.current_state == 5'h04;
  assign _277_ = _275_ | _276_;
  assign _278_ = \rsc0.current_state == 5'h05;
  assign _279_ = _277_ | _278_;
  assign _280_ = \rsc0.current_state == 5'h06;
  assign _281_ = _279_ | _280_;
  assign _282_ = \rsc0.current_state == 5'h07;
  assign _283_ = _281_ | _282_;
  assign _284_ = \rsc0.current_state == 5'h08;
  assign _285_ = _283_ | _284_;
  assign _286_ = \rsc0.current_state == 5'h0f;
  assign _287_ = _285_ | _286_;
  assign _288_ = \rsc0.src_ready & _287_;
  assign _289_ = _274_ | _288_;
  assign _290_ = _289_ ? 1'h1 : 1'h0;
  assign _291_ = \rsc0.src_ready | \rsc0.msg_done ;
  assign _292_ = \rsc0.current_state == 5'h07;
  assign _293_ = \rsc0.current_state == 5'h08;
  assign _294_ = _292_ | _293_;
  assign _295_ = \rsc0.current_state == 5'h05;
  assign _296_ = _294_ | _295_;
  assign _297_ = \rsc0.current_state == 5'h06;
  assign _298_ = _296_ | _297_;
  assign _299_ = \rsc0.current_state == 5'h0e;
  assign _300_ = _298_ | _299_;
  assign _301_ = \rsc0.current_state == 5'h0f;
  assign _302_ = _300_ | _301_;
  assign _303_ = \rsc0.current_state == 5'h0d;
  assign _304_ = _302_ | _303_;
  assign _305_ = _304_ & _291_;
  assign _306_ = \rsc0.current_state == 5'h09;
  assign _307_ = \rsc0.current_state == 5'h0a;
  assign _308_ = _306_ | _307_;
  assign _309_ = \rsc0.current_state == 5'h0b;
  assign _310_ = _308_ | _309_;
  assign _311_ = \rsc0.current_state == 5'h0c;
  assign _312_ = _310_ | _311_;
  assign _313_ = _305_ | _312_;
  assign _314_ = _313_ ? 1'h1 : 1'h0;
  assign _315_ = \rsc0.current_state == 5'h04;
  assign _316_ = \rsc0.current_state == 5'h05;
  assign _317_ = _315_ | _316_;
  assign _318_ = \rsc0.current_state == 5'h06;
  assign _319_ = _317_ | _318_;
  assign _320_ = \rsc0.current_state == 5'h07;
  assign _321_ = _319_ | _320_;
  assign _322_ = \rsc0.current_state == 5'h08;
  assign _323_ = _321_ | _322_;
  assign _324_ = \rsc0.current_state == 5'h0f;
  assign _325_ = _323_ | _324_;
  assign _326_ = _325_ & \rsc0.src_ready ;
  assign _327_ = \rsc0.current_state == 5'h0e;
  assign _328_ = \rsc0.src_ready & _327_;
  assign _329_ = ~\rsc0.msg_done ;
  assign _330_ = _329_ & _328_;
  assign _331_ = _326_ | _330_;
  assign _332_ = \rsc0.current_state == 5'h09;
  assign _333_ = _331_ | _332_;
  assign _334_ = \rsc0.current_state == 5'h0a;
  assign _335_ = _333_ | _334_;
  assign _336_ = \rsc0.current_state == 5'h0b;
  assign _337_ = _335_ | _336_;
  assign _338_ = \rsc0.current_state == 5'h0c;
  assign _339_ = _337_ | _338_;
  assign _340_ = _339_ ? 1'h1 : 1'h0;
  assign _341_ = \rsc0.current_state == 5'h05;
  assign _342_ = \rsc0.current_state == 5'h04;
  assign _343_ = _341_ | _342_;
  assign _344_ = \rsc0.current_state == 5'h06;
  assign _345_ = _343_ | _344_;
  assign _346_ = \rsc0.current_state == 5'h07;
  assign _347_ = _345_ | _346_;
  assign _348_ = \rsc0.current_state == 5'h08;
  assign _349_ = _347_ | _348_;
  assign _350_ = \rsc0.current_state == 5'h0e;
  assign _351_ = \rsc0.current_state == 5'h0f;
  assign _352_ = _350_ | _351_;
  assign _353_ = ~\rsc0.msg_done ;
  assign _354_ = _353_ & _352_;
  assign _355_ = _349_ | _354_;
  assign _356_ = _355_ & \rsc0.src_ready ;
  assign _357_ = \rsc0.current_state == 5'h09;
  assign _358_ = _356_ | _357_;
  assign _359_ = \rsc0.current_state == 5'h0a;
  assign _360_ = _358_ | _359_;
  assign _361_ = \rsc0.current_state == 5'h0b;
  assign _362_ = _360_ | _361_;
  assign _363_ = \rsc0.current_state == 5'h0c;
  assign _364_ = _362_ | _363_;
  assign _365_ = _364_ ? 1'h1 : 1'h0;
  assign _366_ = \rsc0.current_state == 5'h0e;
  assign _367_ = _366_ ? 1'h1 : 1'h0;
  assign _368_ = \rsc0.current_state == 5'h09;
  assign _369_ = \rsc0.current_state == 5'h0a;
  assign _370_ = _368_ | _369_;
  assign _371_ = \rsc0.current_state == 5'h0b;
  assign _372_ = _370_ | _371_;
  assign _373_ = _372_ ? 1'h1 : 1'h0;
  assign _374_ = \rsc0.current_state == 5'h04;
  assign _375_ = \rsc0.current_state == 5'h0e;
  assign _376_ = _374_ | _375_;
  assign _377_ = _376_ ? 1'h1 : 1'h0;
  assign _378_ = \rsc0.current_state == 5'h0e;
  assign _379_ = _378_ ? 1'h1 : 1'h0;
  assign _380_ = \rsc0.current_state == 5'h10;
  assign _381_ = ~\rsc0.dst_ready ;
  assign _382_ = _381_ & _380_;
  assign _383_ = _382_ ? 1'h1 : 1'h0;
  assign _384_ = \rsc0.current_state == 5'h12;
  assign _385_ = _384_ ? 1'h1 : 1'h0;
  assign _386_ = \rsc0.current_state == 5'h11;
  assign _388_ = _386_ ? 1'h1 : 1'h0;
  assign _389_ = \rsc0.current_state == 5'h08;
  assign _390_ = \rsc0.src_ready & _389_;
  assign _391_ = _390_ ? 1'h1 : 1'h0;
  always @(posedge \rsc0.clk , posedge \rsc0.rst )
    if (\rsc0.rst ) _392_ <= 5'h12;
    else _392_ <= \rsc0.next_state ;
  assign _387_ = \rsc0.src_ready ? 5'h01 : 5'h00;
  assign _393_ = !\rsc0.current_state ;
  assign _394_ = \rsc0.src_ready ? 5'h02 : 5'h01;
  assign _395_ = \rsc0.current_state == 5'h01;
  assign _396_ = ~\rsc0.last_block ;
  assign _397_ = _396_ | \rsc0.src_ready ;
  assign _398_ = _397_ ? 5'h03 : 5'h02;
  assign _399_ = \rsc0.current_state == 5'h02;
  assign _400_ = \rsc0.src_ready ? 5'h04 : 5'h03;
  assign _401_ = \rsc0.current_state == 5'h03;
  assign _402_ = \rsc0.src_ready ? 5'h05 : 5'h04;
  assign _403_ = \rsc0.current_state == 5'h04;
  assign _404_ = \rsc0.src_ready ? 5'h06 : 5'h05;
  assign _405_ = \rsc0.current_state == 5'h05;
  assign _406_ = \rsc0.z16 & \rsc0.src_ready ;
  assign _407_ = _406_ ? 5'h07 : 5'h06;
  assign _408_ = \rsc0.current_state == 5'h06;
  assign _409_ = \rsc0.src_ready ? 5'h08 : 5'h07;
  assign _410_ = \rsc0.current_state == 5'h07;
  assign _411_ = \rsc0.src_ready ? 5'h09 : 5'h08;
  assign _412_ = \rsc0.current_state == 5'h08;
  assign _413_ = \rsc0.zlast ? 5'h0a : 5'h09;
  assign z16_reg = _009_;
  assign zlast_reg = _010_;
  assign sel2_reg = _016_;
  assign sel_reg = _017_;
  assign wr_data_reg = _001_;
  assign wr_state_reg = _003_;
  assign wr_len_reg = _005_;
  assign wr_result_reg = _004_;
  assign ctr_ena_reg = _006_;
  assign lb_reg = _014_;
  assign dst_write_reg = _008_;
  assign o8_reg = _012_;
  assign ctrl_rst_reg = _020_;
  assign rst_reg = _011_;
  assign src_ready_reg = _000_;
  assign rst_flags_reg = _022_;
  assign kr_wr_wire = _002_;
  assign wr_chctr_reg = _021_;
  assign msg_done_reg = _015_;
  assign sel_gh_reg = _018_;
  assign sel_gh_reg2 = _019_;
  assign src_read = _007_;
  assign dout = _013_;
  assign dst_write = dst_write_reg;
  assign \rsc0.next_state = _436_;
  assign \rsc0.current_state = _392_;
  assign \rsc0.src_read_sig = _290_;
  assign \rsc0.sel2 = _373_;
  assign \rsc0.sel = _367_;
  assign \rsc0.sel_gh = _377_;
  assign \rsc0.sel_gh2 = _379_;
  assign \rsc0.ctrl_rst = _385_;
  assign \rsc0.wr_chctr = _391_;
  assign \rsc0.rst_flags = _388_;
  assign \rsc0.wr_data = _249_;
  assign \rsc0.kw_wr = _365_;
  assign \rsc0.wr_state = _314_;
  assign \rsc0.wr_result = _261_;
  assign \rsc0.wr_len = _439_;
  assign \rsc0.ctr_ena = _340_;
  assign \rsc0.src_read = \rsc0.src_read_sig ;
  assign \rsc0.dst_write = _383_;
  assign _008_ = \rsc0.dst_write ;
  assign _007_ = \rsc0.src_read ;
  assign _006_ = \rsc0.ctr_ena ;
  assign _005_ = \rsc0.wr_len ;
  assign _004_ = \rsc0.wr_result ;
  assign _003_ = \rsc0.wr_state ;
  assign _002_ = \rsc0.kw_wr ;
  assign _001_ = \rsc0.wr_data ;
  assign _022_ = \rsc0.rst_flags ;
  assign _021_ = \rsc0.wr_chctr ;
  assign _020_ = \rsc0.ctrl_rst ;
  assign _019_ = \rsc0.sel_gh2 ;
  assign _018_ = \rsc0.sel_gh ;
  assign _017_ = \rsc0.sel ;
  assign _016_ = \rsc0.sel2 ;
  assign \rsc0.dst_ready = dst_ready;
  assign \rsc0.src_ready = src_ready_reg;
  assign \rsc0.msg_done = msg_done_reg;
  assign \rsc0.last_block = lb_reg;
  assign \rsc0.o8 = o8_reg;
  assign \rsc0.zlast = zlast_reg;
  assign \rsc0.z16 = z16_reg;
  assign \rsc0.rst = rst;
  assign \rsc0.clk = clk;
  assign \dp256_gen.datapath.from_round = {_037_, _038_, _039_, _040_, _041_, _042_, _043_, _044_};
  assign \dp256_gen.datapath.to_round = {
    \dp256_gen.datapath.st256_gen.sr_gen:1.sr0:438 ,
    \dp256_gen.datapath.st256_gen.sr_gen:2.sr0:442 ,
    \dp256_gen.datapath.st256_gen.sr_gen:3.sr0:446 ,
    \dp256_gen.datapath.st256_gen.sr_gen:4.sr0:450 ,
    \dp256_gen.datapath.st256_gen.sr_gen:5.sr0:454 ,
    \dp256_gen.datapath.st256_gen.sr_gen:6.sr0:458 ,
    \dp256_gen.datapath.st256_gen.sr_gen:7.sr0:462 ,
    \dp256_gen.datapath.st256_gen.sr_gen:8.sr0:466
  };
  assign \dp256_gen.datapath.from_final_add = {
    _045_, \dp256_gen.datapath.result [255:160], _046_, \dp256_gen.datapath.result [127:32]
  };
  assign \dp256_gen.datapath.from_mux = {_047_, _048_, _049_, _050_, _051_, _052_, _053_, _054_};
  assign \dp256_gen.datapath.result = {
    \dp256_gen.datapath.hs256_gen.rr_gen:1.rr:561 ,
    \dp256_gen.datapath.hs256_gen.rr_gen:2.rr:565 ,
    \dp256_gen.datapath.hs256_gen.rr_gen:3.rr:569 ,
    \dp256_gen.datapath.hs256_gen.rr_gen:4.rr:573 ,
    \dp256_gen.datapath.hs256_gen.rr_gen:5.rr:577 ,
    \dp256_gen.datapath.hs256_gen.rr_gen:6.rr:581 ,
    \dp256_gen.datapath.hs256_gen.rr_gen:7.rr:585 ,
    \dp256_gen.datapath.hs256_gen.rr_gen:8.rr:589
  };
  assign \dp256_gen.datapath.to_result = {
    _056_, _057_, _058_, _059_, _060_, _061_, _062_, \dp256_gen.datapath.from_final_add [31:0]
  };
  assign \dp256_gen.datapath.wwire = _071_;
  assign \dp256_gen.datapath.kwire = _078_;
  assign \dp256_gen.datapath.h_exception = _035_;
  assign \dp256_gen.datapath.rd_num = _072_;
  assign \dp256_gen.datapath.z16_reg = _074_;
  assign \dp256_gen.datapath.ena_reg = _055_;
  assign \dp256_gen.datapath.kwhwire = _036_;
  assign \dp256_gen.datapath.kwhreg = \dp256_gen.datapath.kwh_reg:469 ;
  assign \dp256_gen.datapath.chunk_ctr = \dp256_gen.datapath.decounter_gen:603 ;
  assign \dp256_gen.datapath.out_ctr = _077_;
  assign \dp256_gen.datapath.gh = {\dp256_gen.datapath.sel_gh , \dp256_gen.datapath.sel_gh2 };
  assign \dp256_gen.datapath.last_block_out = _073_;
  assign \dp256_gen.datapath.st256_gen.sr_gen:1.sr0:438 = _023_;
  assign \dp256_gen.datapath.st256_gen.sr_gen:2.sr0:442 = _024_;
  assign \dp256_gen.datapath.st256_gen.sr_gen:3.sr0:446 = _025_;
  assign \dp256_gen.datapath.st256_gen.sr_gen:4.sr0:450 = _026_;
  assign \dp256_gen.datapath.st256_gen.sr_gen:5.sr0:454 = _027_;
  assign \dp256_gen.datapath.st256_gen.sr_gen:6.sr0:458 = _028_;
  assign \dp256_gen.datapath.st256_gen.sr_gen:7.sr0:462 = _029_;
  assign \dp256_gen.datapath.st256_gen.sr_gen:8.sr0:466 = _030_;
  assign \dp256_gen.datapath.kwh_reg:469 = _031_;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:1.rr:561 = _063_;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:2.rr:565 = _064_;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:3.rr:569 = _065_;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:4.rr:573 = _066_;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:5.rr:577 = _067_;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:6.rr:581 = _068_;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:7.rr:585 = _069_;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:8.rr:589 = _070_;
  assign \dp256_gen.datapath.decounter_gen:603 = _079_;
  assign \dp256_gen.datapath.z16 = \dp256_gen.datapath.z16_reg ;
  assign \dp256_gen.datapath.zlast = _075_;
  assign \dp256_gen.datapath.o8 = _076_;
  assign \dp256_gen.datapath.dataout = \dp256_gen.datapath.result [255:224];
  assign \dp256_gen.datapath.last_block = \dp256_gen.datapath.last_block_out ;
  assign \dp256_gen.datapath.msg_done = _081_;
  assign \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.output = _225_;
  assign _023_ = \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.output ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.input = \dp256_gen.datapath.from_mux [255:224];
  assign \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.en = \dp256_gen.datapath.wr_state ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:1.sr0.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.output = _228_;
  assign _024_ = \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.output ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.input = \dp256_gen.datapath.from_mux [223:192];
  assign \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.en = \dp256_gen.datapath.wr_state ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:2.sr0.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.output = _231_;
  assign _025_ = \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.output ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.input = \dp256_gen.datapath.from_mux [191:160];
  assign \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.en = \dp256_gen.datapath.wr_state ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:3.sr0.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.output = _234_;
  assign _026_ = \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.output ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.input = \dp256_gen.datapath.from_mux [159:128];
  assign \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.en = \dp256_gen.datapath.wr_state ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:4.sr0.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.output = _237_;
  assign _027_ = \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.output ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.input = \dp256_gen.datapath.from_mux [127:96];
  assign \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.en = \dp256_gen.datapath.wr_state ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:5.sr0.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.output = _240_;
  assign _028_ = \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.output ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.input = \dp256_gen.datapath.from_mux [95:64];
  assign \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.en = \dp256_gen.datapath.wr_state ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:6.sr0.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.output = _243_;
  assign _029_ = \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.output ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.input = \dp256_gen.datapath.from_mux [63:32];
  assign \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.en = \dp256_gen.datapath.wr_state ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:7.sr0.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.output = _246_;
  assign _030_ = \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.output ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.input = \dp256_gen.datapath.from_mux [31:0];
  assign \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.en = \dp256_gen.datapath.wr_state ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.st256_gen.sr_gen:8.sr0.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.kwh_reg.output = _185_;
  assign _031_ = \dp256_gen.datapath.kwh_reg.output ;
  assign \dp256_gen.datapath.kwh_reg.input = \dp256_gen.datapath.kwhwire ;
  assign \dp256_gen.datapath.kwh_reg.en = \dp256_gen.datapath.kw_wr ;
  assign \dp256_gen.datapath.kwh_reg.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.kwh_reg.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.round.cf0_reg = _196_;
  assign \dp256_gen.datapath.round.cf1_reg = _197_;
  assign \dp256_gen.datapath.round.ch_reg = _198_;
  assign \dp256_gen.datapath.round.maj_reg = _199_;
  assign \dp256_gen.datapath.round.g_or_h = _207_;
  assign \dp256_gen.datapath.round.kwhwire = _209_;
  assign \dp256_gen.datapath.round.aout = _206_;
  assign \dp256_gen.datapath.round.bout = \dp256_gen.datapath.round.ain ;
  assign \dp256_gen.datapath.round.cout = \dp256_gen.datapath.round.bin ;
  assign \dp256_gen.datapath.round.dout = \dp256_gen.datapath.round.cin ;
  assign \dp256_gen.datapath.round.eout = _202_;
  assign \dp256_gen.datapath.round.fout = \dp256_gen.datapath.round.ein ;
  assign \dp256_gen.datapath.round.gout = \dp256_gen.datapath.round.fin ;
  assign \dp256_gen.datapath.round.hout = \dp256_gen.datapath.round.gin ;
  assign \dp256_gen.datapath.round.a32.s0.tmp = \dp256_gen.datapath.round.a32.s0.x [21:0];
  assign \dp256_gen.datapath.round.a32.s0.o = _211_;
  assign _196_ = \dp256_gen.datapath.round.a32.s0.o ;
  assign \dp256_gen.datapath.round.a32.s0.x = \dp256_gen.datapath.round.ain ;
  assign \dp256_gen.datapath.round.a32.s1.tmp = \dp256_gen.datapath.round.a32.s1.x [24:0];
  assign \dp256_gen.datapath.round.a32.s1.o = _213_;
  assign _197_ = \dp256_gen.datapath.round.a32.s1.o ;
  assign \dp256_gen.datapath.round.a32.s1.x = \dp256_gen.datapath.round.ein ;
  assign \dp256_gen.datapath.round.c1.o = _217_;
  assign _198_ = \dp256_gen.datapath.round.c1.o ;
  assign \dp256_gen.datapath.round.c1.z = \dp256_gen.datapath.round.gin ;
  assign \dp256_gen.datapath.round.c1.y = \dp256_gen.datapath.round.fin ;
  assign \dp256_gen.datapath.round.c1.x = \dp256_gen.datapath.round.ein ;
  assign \dp256_gen.datapath.round.m1.o = _222_;
  assign _199_ = \dp256_gen.datapath.round.m1.o ;
  assign \dp256_gen.datapath.round.m1.z = \dp256_gen.datapath.round.cin ;
  assign \dp256_gen.datapath.round.m1.y = \dp256_gen.datapath.round.bin ;
  assign \dp256_gen.datapath.round.m1.x = \dp256_gen.datapath.round.ain ;
  assign _044_ = \dp256_gen.datapath.round.hout ;
  assign _043_ = \dp256_gen.datapath.round.gout ;
  assign _042_ = \dp256_gen.datapath.round.fout ;
  assign _041_ = \dp256_gen.datapath.round.eout ;
  assign _040_ = \dp256_gen.datapath.round.dout ;
  assign _039_ = \dp256_gen.datapath.round.cout ;
  assign _038_ = \dp256_gen.datapath.round.bout ;
  assign _037_ = \dp256_gen.datapath.round.aout ;
  assign _036_ = \dp256_gen.datapath.round.kwhwire ;
  assign \dp256_gen.datapath.round.hin = \dp256_gen.datapath.h_exception ;
  assign \dp256_gen.datapath.round.gin = \dp256_gen.datapath.to_round [63:32];
  assign \dp256_gen.datapath.round.fin = \dp256_gen.datapath.to_round [95:64];
  assign \dp256_gen.datapath.round.ein = \dp256_gen.datapath.to_round [127:96];
  assign \dp256_gen.datapath.round.din = \dp256_gen.datapath.to_round [159:128];
  assign \dp256_gen.datapath.round.cin = \dp256_gen.datapath.to_round [191:160];
  assign \dp256_gen.datapath.round.bin = \dp256_gen.datapath.to_round [223:192];
  assign \dp256_gen.datapath.round.ain = \dp256_gen.datapath.to_round [255:224];
  assign \dp256_gen.datapath.round.wwire = \dp256_gen.datapath.wwire ;
  assign \dp256_gen.datapath.round.kwire = \dp256_gen.datapath.kwire ;
  assign \dp256_gen.datapath.round.kw = \dp256_gen.datapath.kwhreg ;
  assign \dp256_gen.datapath.round.sel_gh = \dp256_gen.datapath.sel_gh ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.output = _161_;
  assign _063_ = \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.output ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.input = \dp256_gen.datapath.to_result [255:224];
  assign \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.en = \dp256_gen.datapath.ena_reg ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:1.rr.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.output = _164_;
  assign _064_ = \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.output ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.input = \dp256_gen.datapath.to_result [223:192];
  assign \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.en = \dp256_gen.datapath.ena_reg ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:2.rr.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.output = _167_;
  assign _065_ = \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.output ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.input = \dp256_gen.datapath.to_result [191:160];
  assign \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.en = \dp256_gen.datapath.ena_reg ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:3.rr.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.output = _170_;
  assign _066_ = \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.output ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.input = \dp256_gen.datapath.to_result [159:128];
  assign \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.en = \dp256_gen.datapath.ena_reg ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:4.rr.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.output = _173_;
  assign _067_ = \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.output ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.input = \dp256_gen.datapath.to_result [127:96];
  assign \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.en = \dp256_gen.datapath.ena_reg ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:5.rr.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.output = _176_;
  assign _068_ = \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.output ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.input = \dp256_gen.datapath.to_result [95:64];
  assign \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.en = \dp256_gen.datapath.ena_reg ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:6.rr.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.output = _179_;
  assign _069_ = \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.output ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.input = \dp256_gen.datapath.to_result [63:32];
  assign \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.en = \dp256_gen.datapath.ena_reg ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:7.rr.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.output = _182_;
  assign _070_ = \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.output ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.input = \dp256_gen.datapath.to_result [31:0];
  assign \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.en = \dp256_gen.datapath.ena_reg ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.hs256_gen.rr_gen:8.rr.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.dc.wires = {
    _103_,
    _142_,
    _140_,
    _138_,
    _136_,
    _134_,
    _132_,
    _130_,
    _128_,
    _126_,
    _124_,
    _122_,
    _120_,
    _118_,
    _116_,
    _114_,
    _112_
  };
  assign \dp256_gen.datapath.dc.wwires = _110_;
  assign \dp256_gen.datapath.dc.d_one_wire = _105_;
  assign \dp256_gen.datapath.dc.d_zero_wire = _104_;
  assign \dp256_gen.datapath.dc.first_stage = _106_;
  assign \dp256_gen.datapath.dc.to_second_stage = _107_;
  assign \dp256_gen.datapath.dc.second_stage = _108_;
  assign \dp256_gen.datapath.dc.to_third_stage = _109_;
  assign \dp256_gen.datapath.dc.w = \dp256_gen.datapath.dc.wires [511:480];
  assign \dp256_gen.datapath.dc.a32.d0.tmp = 3'h0;
  assign \dp256_gen.datapath.dc.a32.d0.o = _144_;
  assign _104_ = \dp256_gen.datapath.dc.a32.d0.o ;
  assign \dp256_gen.datapath.dc.a32.d0.x = \dp256_gen.datapath.dc.wires [127:96];
  assign \dp256_gen.datapath.dc.a32.d1.tmp = 10'h000;
  assign \dp256_gen.datapath.dc.a32.d1.o = _146_;
  assign _105_ = \dp256_gen.datapath.dc.a32.d1.o ;
  assign \dp256_gen.datapath.dc.a32.d1.x = \dp256_gen.datapath.dc.wires [479:448];
  assign \dp256_gen.datapath.dc.reg01.output = _149_;
  assign _107_ = \dp256_gen.datapath.dc.reg01.output ;
  assign \dp256_gen.datapath.dc.reg01.input = \dp256_gen.datapath.dc.first_stage ;
  assign \dp256_gen.datapath.dc.reg01.en = \dp256_gen.datapath.dc.wr_data ;
  assign \dp256_gen.datapath.dc.reg01.rst = 1'h0;
  assign \dp256_gen.datapath.dc.reg01.clk = \dp256_gen.datapath.dc.clk ;
  assign \dp256_gen.datapath.dc.reg02.output = _152_;
  assign _109_ = \dp256_gen.datapath.dc.reg02.output ;
  assign \dp256_gen.datapath.dc.reg02.input = \dp256_gen.datapath.dc.second_stage ;
  assign \dp256_gen.datapath.dc.reg02.en = \dp256_gen.datapath.dc.wr_data ;
  assign \dp256_gen.datapath.dc.reg02.rst = 1'h0;
  assign \dp256_gen.datapath.dc.reg02.clk = \dp256_gen.datapath.dc.clk ;
  assign _071_ = \dp256_gen.datapath.dc.w ;
  assign \dp256_gen.datapath.dc.data = \dp256_gen.datapath.data ;
  assign \dp256_gen.datapath.dc.wr_data = \dp256_gen.datapath.wr_data ;
  assign \dp256_gen.datapath.dc.sel = \dp256_gen.datapath.sel2 ;
  assign \dp256_gen.datapath.dc.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.rd_ctr.reg = _195_;
  assign \dp256_gen.datapath.rd_ctr.ctr = \dp256_gen.datapath.rd_ctr.reg ;
  assign _072_ = \dp256_gen.datapath.rd_ctr.ctr ;
  assign \dp256_gen.datapath.rd_ctr.ena = \dp256_gen.datapath.ctr_ena ;
  assign \dp256_gen.datapath.rd_ctr.reset = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.rd_ctr.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.bf.z16_in = _083_;
  assign \dp256_gen.datapath.bf.z16_out = \dp256_gen.datapath.bf.r0:979 ;
  assign \dp256_gen.datapath.bf.zlast_in = _085_;
  assign \dp256_gen.datapath.bf.zlast_out = \dp256_gen.datapath.bf.r1:982 ;
  assign \dp256_gen.datapath.bf.o8_in = _087_;
  assign \dp256_gen.datapath.bf.r0:979 = _088_;
  assign \dp256_gen.datapath.bf.r1:982 = _089_;
  assign \dp256_gen.datapath.bf.r4:985 = _090_;
  assign \dp256_gen.datapath.bf.last_block_out = \dp256_gen.datapath.bf.r4:985 ;
  assign \dp256_gen.datapath.bf.z16 = \dp256_gen.datapath.bf.z16_out ;
  assign \dp256_gen.datapath.bf.zlast = \dp256_gen.datapath.bf.zlast_out ;
  assign \dp256_gen.datapath.bf.o8 = \dp256_gen.datapath.bf.o8_in ;
  assign \dp256_gen.datapath.bf.r0.r = _093_;
  assign \dp256_gen.datapath.bf.r0.q = \dp256_gen.datapath.bf.r0.r ;
  assign _088_ = \dp256_gen.datapath.bf.r0.q ;
  assign \dp256_gen.datapath.bf.r0.d = \dp256_gen.datapath.bf.z16_in ;
  assign \dp256_gen.datapath.bf.r0.rst = \dp256_gen.datapath.bf.rst ;
  assign \dp256_gen.datapath.bf.r0.ena = \dp256_gen.datapath.bf.en ;
  assign \dp256_gen.datapath.bf.r0.clk = \dp256_gen.datapath.bf.clk ;
  assign \dp256_gen.datapath.bf.r1.r = _096_;
  assign \dp256_gen.datapath.bf.r1.q = \dp256_gen.datapath.bf.r1.r ;
  assign _089_ = \dp256_gen.datapath.bf.r1.q ;
  assign \dp256_gen.datapath.bf.r1.d = \dp256_gen.datapath.bf.zlast_in ;
  assign \dp256_gen.datapath.bf.r1.rst = \dp256_gen.datapath.bf.rst ;
  assign \dp256_gen.datapath.bf.r1.ena = \dp256_gen.datapath.bf.en ;
  assign \dp256_gen.datapath.bf.r1.clk = \dp256_gen.datapath.bf.clk ;
  assign \dp256_gen.datapath.bf.r4.r = _099_;
  assign \dp256_gen.datapath.bf.r4.q = \dp256_gen.datapath.bf.r4.r ;
  assign _090_ = \dp256_gen.datapath.bf.r4.q ;
  assign \dp256_gen.datapath.bf.r4.d = \dp256_gen.datapath.bf.last_block_in ;
  assign \dp256_gen.datapath.bf.r4.rst = \dp256_gen.datapath.bf.rst_flags ;
  assign \dp256_gen.datapath.bf.r4.ena = \dp256_gen.datapath.bf.wr_len ;
  assign \dp256_gen.datapath.bf.r4.clk = \dp256_gen.datapath.bf.clk ;
  assign _076_ = \dp256_gen.datapath.bf.o8 ;
  assign _075_ = \dp256_gen.datapath.bf.zlast ;
  assign _074_ = \dp256_gen.datapath.bf.z16 ;
  assign _073_ = \dp256_gen.datapath.bf.last_block_out ;
  assign \dp256_gen.datapath.bf.rst_flags = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.bf.rst = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.bf.out_ctr = \dp256_gen.datapath.out_ctr ;
  assign \dp256_gen.datapath.bf.exam_block = \dp256_gen.datapath.data ;
  assign \dp256_gen.datapath.bf.rd_num = \dp256_gen.datapath.rd_num ;
  assign \dp256_gen.datapath.bf.last_block_in = \dp256_gen.datapath.data [31];
  assign \dp256_gen.datapath.bf.wr_len = \dp256_gen.datapath.wr_len ;
  assign \dp256_gen.datapath.bf.en = \dp256_gen.datapath.ctr_ena ;
  assign \dp256_gen.datapath.bf.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.o_ctr.reg = _190_;
  assign \dp256_gen.datapath.o_ctr.ctr = \dp256_gen.datapath.o_ctr.reg ;
  assign _077_ = \dp256_gen.datapath.o_ctr.ctr ;
  assign \dp256_gen.datapath.o_ctr.ena = \dp256_gen.datapath.dst_write ;
  assign \dp256_gen.datapath.o_ctr.reset = \dp256_gen.datapath.rst ;
  assign \dp256_gen.datapath.o_ctr.clk = \dp256_gen.datapath.clk ;
  assign \dp256_gen.datapath.const.output = _102_;
  assign _078_ = \dp256_gen.datapath.const.output ;
  assign \dp256_gen.datapath.const.address = \dp256_gen.datapath.rd_num ;
  assign \dp256_gen.datapath.decounter_gen.reg_in = _153_;
  assign \dp256_gen.datapath.decounter_gen.reg_out = _158_;
  assign \dp256_gen.datapath.decounter_gen.ctrl = _155_;
  assign \dp256_gen.datapath.decounter_gen.output = \dp256_gen.datapath.decounter_gen.reg_out ;
  assign _079_ = \dp256_gen.datapath.decounter_gen.output ;
  assign \dp256_gen.datapath.decounter_gen.input = \dp256_gen.datapath.data [30:9];
  assign \dp256_gen.datapath.decounter_gen.en = \dp256_gen.datapath.wr_chctr ;
  assign \dp256_gen.datapath.decounter_gen.load = \dp256_gen.datapath.wr_len ;
  assign \dp256_gen.datapath.decounter_gen.rst = 1'h0;
  assign \dp256_gen.datapath.decounter_gen.clk = \dp256_gen.datapath.clk ;
  assign _015_ = \dp256_gen.datapath.msg_done ;
  assign _014_ = \dp256_gen.datapath.last_block ;
  assign _013_ = \dp256_gen.datapath.dataout ;
  assign _012_ = \dp256_gen.datapath.o8 ;
  assign _010_ = \dp256_gen.datapath.zlast ;
  assign _009_ = \dp256_gen.datapath.z16 ;
  assign \dp256_gen.datapath.rst_flags = rst_flags_reg;
  assign \dp256_gen.datapath.wr_chctr = wr_chctr_reg;
  assign \dp256_gen.datapath.data = din;
  assign \dp256_gen.datapath.dst_write = dst_write_reg;
  assign \dp256_gen.datapath.ctr_ena = ctr_ena_reg;
  assign \dp256_gen.datapath.sel_gh2 = sel_gh_reg2;
  assign \dp256_gen.datapath.sel_gh = sel_gh_reg;
  assign \dp256_gen.datapath.sel2 = sel2_reg;
  assign \dp256_gen.datapath.sel = sel_reg;
  assign \dp256_gen.datapath.wr_len = wr_len_reg;
  assign \dp256_gen.datapath.kw_wr = kr_wr_wire;
  assign \dp256_gen.datapath.wr_data = wr_data_reg;
  assign \dp256_gen.datapath.wr_result = wr_result_reg;
  assign \dp256_gen.datapath.wr_state = wr_state_reg;
  assign \dp256_gen.datapath.rst = rst_reg;
  assign \dp256_gen.datapath.clk = clk;
endmodule
