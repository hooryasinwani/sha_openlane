module sha2_top (clk,
    dst_ready,
    dst_write,
    rst,
    src_read,
    src_ready,
    din,
    dout);
 input clk;
 input dst_ready;
 output dst_write;
 input rst;
 output src_read;
 input src_ready;
 input [31:0] din;
 output [31:0] dout;

 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _093_;
 wire _096_;
 wire _099_;
 wire \_116_[0] ;
 wire \_116_[10] ;
 wire \_116_[11] ;
 wire \_116_[12] ;
 wire \_116_[13] ;
 wire \_116_[14] ;
 wire \_116_[15] ;
 wire \_116_[16] ;
 wire \_116_[17] ;
 wire \_116_[18] ;
 wire \_116_[19] ;
 wire \_116_[1] ;
 wire \_116_[20] ;
 wire \_116_[21] ;
 wire \_116_[22] ;
 wire \_116_[23] ;
 wire \_116_[24] ;
 wire \_116_[25] ;
 wire \_116_[26] ;
 wire \_116_[27] ;
 wire \_116_[28] ;
 wire \_116_[29] ;
 wire \_116_[2] ;
 wire \_116_[30] ;
 wire \_116_[31] ;
 wire \_116_[3] ;
 wire \_116_[4] ;
 wire \_116_[5] ;
 wire \_116_[6] ;
 wire \_116_[7] ;
 wire \_116_[8] ;
 wire \_116_[9] ;
 wire \_118_[0] ;
 wire \_118_[10] ;
 wire \_118_[11] ;
 wire \_118_[12] ;
 wire \_118_[13] ;
 wire \_118_[14] ;
 wire \_118_[15] ;
 wire \_118_[16] ;
 wire \_118_[17] ;
 wire \_118_[18] ;
 wire \_118_[19] ;
 wire \_118_[1] ;
 wire \_118_[20] ;
 wire \_118_[21] ;
 wire \_118_[22] ;
 wire \_118_[23] ;
 wire \_118_[24] ;
 wire \_118_[25] ;
 wire \_118_[26] ;
 wire \_118_[27] ;
 wire \_118_[28] ;
 wire \_118_[29] ;
 wire \_118_[2] ;
 wire \_118_[30] ;
 wire \_118_[31] ;
 wire \_118_[3] ;
 wire \_118_[4] ;
 wire \_118_[5] ;
 wire \_118_[6] ;
 wire \_118_[7] ;
 wire \_118_[8] ;
 wire \_118_[9] ;
 wire \_120_[0] ;
 wire \_120_[10] ;
 wire \_120_[11] ;
 wire \_120_[12] ;
 wire \_120_[13] ;
 wire \_120_[14] ;
 wire \_120_[15] ;
 wire \_120_[16] ;
 wire \_120_[17] ;
 wire \_120_[18] ;
 wire \_120_[19] ;
 wire \_120_[1] ;
 wire \_120_[20] ;
 wire \_120_[21] ;
 wire \_120_[22] ;
 wire \_120_[23] ;
 wire \_120_[24] ;
 wire \_120_[25] ;
 wire \_120_[26] ;
 wire \_120_[27] ;
 wire \_120_[28] ;
 wire \_120_[29] ;
 wire \_120_[2] ;
 wire \_120_[30] ;
 wire \_120_[31] ;
 wire \_120_[3] ;
 wire \_120_[4] ;
 wire \_120_[5] ;
 wire \_120_[6] ;
 wire \_120_[7] ;
 wire \_120_[8] ;
 wire \_120_[9] ;
 wire \_122_[0] ;
 wire \_122_[10] ;
 wire \_122_[11] ;
 wire \_122_[12] ;
 wire \_122_[13] ;
 wire \_122_[14] ;
 wire \_122_[15] ;
 wire \_122_[16] ;
 wire \_122_[17] ;
 wire \_122_[18] ;
 wire \_122_[19] ;
 wire \_122_[1] ;
 wire \_122_[20] ;
 wire \_122_[21] ;
 wire \_122_[22] ;
 wire \_122_[23] ;
 wire \_122_[24] ;
 wire \_122_[25] ;
 wire \_122_[26] ;
 wire \_122_[27] ;
 wire \_122_[28] ;
 wire \_122_[29] ;
 wire \_122_[2] ;
 wire \_122_[30] ;
 wire \_122_[31] ;
 wire \_122_[3] ;
 wire \_122_[4] ;
 wire \_122_[5] ;
 wire \_122_[6] ;
 wire \_122_[7] ;
 wire \_122_[8] ;
 wire \_122_[9] ;
 wire \_124_[0] ;
 wire \_124_[10] ;
 wire \_124_[11] ;
 wire \_124_[12] ;
 wire \_124_[13] ;
 wire \_124_[14] ;
 wire \_124_[15] ;
 wire \_124_[16] ;
 wire \_124_[17] ;
 wire \_124_[18] ;
 wire \_124_[19] ;
 wire \_124_[1] ;
 wire \_124_[20] ;
 wire \_124_[21] ;
 wire \_124_[22] ;
 wire \_124_[23] ;
 wire \_124_[24] ;
 wire \_124_[25] ;
 wire \_124_[26] ;
 wire \_124_[27] ;
 wire \_124_[28] ;
 wire \_124_[29] ;
 wire \_124_[2] ;
 wire \_124_[30] ;
 wire \_124_[31] ;
 wire \_124_[3] ;
 wire \_124_[4] ;
 wire \_124_[5] ;
 wire \_124_[6] ;
 wire \_124_[7] ;
 wire \_124_[8] ;
 wire \_124_[9] ;
 wire \_126_[0] ;
 wire \_126_[10] ;
 wire \_126_[11] ;
 wire \_126_[12] ;
 wire \_126_[13] ;
 wire \_126_[14] ;
 wire \_126_[15] ;
 wire \_126_[16] ;
 wire \_126_[17] ;
 wire \_126_[18] ;
 wire \_126_[19] ;
 wire \_126_[1] ;
 wire \_126_[20] ;
 wire \_126_[21] ;
 wire \_126_[22] ;
 wire \_126_[23] ;
 wire \_126_[24] ;
 wire \_126_[25] ;
 wire \_126_[26] ;
 wire \_126_[27] ;
 wire \_126_[28] ;
 wire \_126_[29] ;
 wire \_126_[2] ;
 wire \_126_[30] ;
 wire \_126_[31] ;
 wire \_126_[3] ;
 wire \_126_[4] ;
 wire \_126_[5] ;
 wire \_126_[6] ;
 wire \_126_[7] ;
 wire \_126_[8] ;
 wire \_126_[9] ;
 wire \_128_[0] ;
 wire \_128_[10] ;
 wire \_128_[11] ;
 wire \_128_[12] ;
 wire \_128_[13] ;
 wire \_128_[14] ;
 wire \_128_[15] ;
 wire \_128_[16] ;
 wire \_128_[17] ;
 wire \_128_[18] ;
 wire \_128_[19] ;
 wire \_128_[1] ;
 wire \_128_[20] ;
 wire \_128_[21] ;
 wire \_128_[22] ;
 wire \_128_[23] ;
 wire \_128_[24] ;
 wire \_128_[25] ;
 wire \_128_[26] ;
 wire \_128_[27] ;
 wire \_128_[28] ;
 wire \_128_[29] ;
 wire \_128_[2] ;
 wire \_128_[30] ;
 wire \_128_[31] ;
 wire \_128_[3] ;
 wire \_128_[4] ;
 wire \_128_[5] ;
 wire \_128_[6] ;
 wire \_128_[7] ;
 wire \_128_[8] ;
 wire \_128_[9] ;
 wire \_130_[0] ;
 wire \_130_[10] ;
 wire \_130_[11] ;
 wire \_130_[12] ;
 wire \_130_[13] ;
 wire \_130_[14] ;
 wire \_130_[15] ;
 wire \_130_[16] ;
 wire \_130_[17] ;
 wire \_130_[18] ;
 wire \_130_[19] ;
 wire \_130_[1] ;
 wire \_130_[20] ;
 wire \_130_[21] ;
 wire \_130_[22] ;
 wire \_130_[23] ;
 wire \_130_[24] ;
 wire \_130_[25] ;
 wire \_130_[26] ;
 wire \_130_[27] ;
 wire \_130_[28] ;
 wire \_130_[29] ;
 wire \_130_[2] ;
 wire \_130_[30] ;
 wire \_130_[31] ;
 wire \_130_[3] ;
 wire \_130_[4] ;
 wire \_130_[5] ;
 wire \_130_[6] ;
 wire \_130_[7] ;
 wire \_130_[8] ;
 wire \_130_[9] ;
 wire \_132_[0] ;
 wire \_132_[10] ;
 wire \_132_[11] ;
 wire \_132_[12] ;
 wire \_132_[13] ;
 wire \_132_[14] ;
 wire \_132_[15] ;
 wire \_132_[16] ;
 wire \_132_[17] ;
 wire \_132_[18] ;
 wire \_132_[19] ;
 wire \_132_[1] ;
 wire \_132_[20] ;
 wire \_132_[21] ;
 wire \_132_[22] ;
 wire \_132_[23] ;
 wire \_132_[24] ;
 wire \_132_[25] ;
 wire \_132_[26] ;
 wire \_132_[27] ;
 wire \_132_[28] ;
 wire \_132_[29] ;
 wire \_132_[2] ;
 wire \_132_[30] ;
 wire \_132_[31] ;
 wire \_132_[3] ;
 wire \_132_[4] ;
 wire \_132_[5] ;
 wire \_132_[6] ;
 wire \_132_[7] ;
 wire \_132_[8] ;
 wire \_132_[9] ;
 wire \_134_[0] ;
 wire \_134_[10] ;
 wire \_134_[11] ;
 wire \_134_[12] ;
 wire \_134_[13] ;
 wire \_134_[14] ;
 wire \_134_[15] ;
 wire \_134_[16] ;
 wire \_134_[17] ;
 wire \_134_[18] ;
 wire \_134_[19] ;
 wire \_134_[1] ;
 wire \_134_[20] ;
 wire \_134_[21] ;
 wire \_134_[22] ;
 wire \_134_[23] ;
 wire \_134_[24] ;
 wire \_134_[25] ;
 wire \_134_[26] ;
 wire \_134_[27] ;
 wire \_134_[28] ;
 wire \_134_[29] ;
 wire \_134_[2] ;
 wire \_134_[30] ;
 wire \_134_[31] ;
 wire \_134_[3] ;
 wire \_134_[4] ;
 wire \_134_[5] ;
 wire \_134_[6] ;
 wire \_134_[7] ;
 wire \_134_[8] ;
 wire \_134_[9] ;
 wire \_136_[0] ;
 wire \_136_[10] ;
 wire \_136_[11] ;
 wire \_136_[12] ;
 wire \_136_[13] ;
 wire \_136_[14] ;
 wire \_136_[15] ;
 wire \_136_[16] ;
 wire \_136_[17] ;
 wire \_136_[18] ;
 wire \_136_[19] ;
 wire \_136_[1] ;
 wire \_136_[20] ;
 wire \_136_[21] ;
 wire \_136_[22] ;
 wire \_136_[23] ;
 wire \_136_[24] ;
 wire \_136_[25] ;
 wire \_136_[26] ;
 wire \_136_[27] ;
 wire \_136_[28] ;
 wire \_136_[29] ;
 wire \_136_[2] ;
 wire \_136_[30] ;
 wire \_136_[31] ;
 wire \_136_[3] ;
 wire \_136_[4] ;
 wire \_136_[5] ;
 wire \_136_[6] ;
 wire \_136_[7] ;
 wire \_136_[8] ;
 wire \_136_[9] ;
 wire \_138_[0] ;
 wire \_138_[10] ;
 wire \_138_[11] ;
 wire \_138_[12] ;
 wire \_138_[13] ;
 wire \_138_[14] ;
 wire \_138_[15] ;
 wire \_138_[16] ;
 wire \_138_[17] ;
 wire \_138_[18] ;
 wire \_138_[19] ;
 wire \_138_[1] ;
 wire \_138_[20] ;
 wire \_138_[21] ;
 wire \_138_[22] ;
 wire \_138_[23] ;
 wire \_138_[24] ;
 wire \_138_[25] ;
 wire \_138_[26] ;
 wire \_138_[27] ;
 wire \_138_[28] ;
 wire \_138_[29] ;
 wire \_138_[2] ;
 wire \_138_[30] ;
 wire \_138_[31] ;
 wire \_138_[3] ;
 wire \_138_[4] ;
 wire \_138_[5] ;
 wire \_138_[6] ;
 wire \_138_[7] ;
 wire \_138_[8] ;
 wire \_138_[9] ;
 wire \_140_[0] ;
 wire \_140_[10] ;
 wire \_140_[11] ;
 wire \_140_[12] ;
 wire \_140_[13] ;
 wire \_140_[14] ;
 wire \_140_[15] ;
 wire \_140_[16] ;
 wire \_140_[17] ;
 wire \_140_[18] ;
 wire \_140_[19] ;
 wire \_140_[1] ;
 wire \_140_[20] ;
 wire \_140_[21] ;
 wire \_140_[22] ;
 wire \_140_[23] ;
 wire \_140_[24] ;
 wire \_140_[25] ;
 wire \_140_[26] ;
 wire \_140_[27] ;
 wire \_140_[28] ;
 wire \_140_[29] ;
 wire \_140_[2] ;
 wire \_140_[30] ;
 wire \_140_[31] ;
 wire \_140_[3] ;
 wire \_140_[4] ;
 wire \_140_[5] ;
 wire \_140_[6] ;
 wire \_140_[7] ;
 wire \_140_[8] ;
 wire \_140_[9] ;
 wire \_142_[0] ;
 wire \_142_[10] ;
 wire \_142_[11] ;
 wire \_142_[12] ;
 wire \_142_[13] ;
 wire \_142_[14] ;
 wire \_142_[15] ;
 wire \_142_[16] ;
 wire \_142_[17] ;
 wire \_142_[18] ;
 wire \_142_[19] ;
 wire \_142_[1] ;
 wire \_142_[20] ;
 wire \_142_[21] ;
 wire \_142_[22] ;
 wire \_142_[23] ;
 wire \_142_[24] ;
 wire \_142_[25] ;
 wire \_142_[26] ;
 wire \_142_[27] ;
 wire \_142_[28] ;
 wire \_142_[29] ;
 wire \_142_[2] ;
 wire \_142_[30] ;
 wire \_142_[31] ;
 wire \_142_[3] ;
 wire \_142_[4] ;
 wire \_142_[5] ;
 wire \_142_[6] ;
 wire \_142_[7] ;
 wire \_142_[8] ;
 wire \_142_[9] ;
 wire \_149_[0] ;
 wire \_149_[10] ;
 wire \_149_[11] ;
 wire \_149_[12] ;
 wire \_149_[13] ;
 wire \_149_[14] ;
 wire \_149_[15] ;
 wire \_149_[16] ;
 wire \_149_[17] ;
 wire \_149_[18] ;
 wire \_149_[19] ;
 wire \_149_[1] ;
 wire \_149_[20] ;
 wire \_149_[21] ;
 wire \_149_[22] ;
 wire \_149_[23] ;
 wire \_149_[24] ;
 wire \_149_[25] ;
 wire \_149_[26] ;
 wire \_149_[27] ;
 wire \_149_[28] ;
 wire \_149_[29] ;
 wire \_149_[2] ;
 wire \_149_[30] ;
 wire \_149_[31] ;
 wire \_149_[3] ;
 wire \_149_[4] ;
 wire \_149_[5] ;
 wire \_149_[6] ;
 wire \_149_[7] ;
 wire \_149_[8] ;
 wire \_149_[9] ;
 wire \_152_[0] ;
 wire \_152_[10] ;
 wire \_152_[11] ;
 wire \_152_[12] ;
 wire \_152_[13] ;
 wire \_152_[14] ;
 wire \_152_[15] ;
 wire \_152_[16] ;
 wire \_152_[17] ;
 wire \_152_[18] ;
 wire \_152_[19] ;
 wire \_152_[1] ;
 wire \_152_[20] ;
 wire \_152_[21] ;
 wire \_152_[22] ;
 wire \_152_[23] ;
 wire \_152_[24] ;
 wire \_152_[25] ;
 wire \_152_[26] ;
 wire \_152_[27] ;
 wire \_152_[28] ;
 wire \_152_[29] ;
 wire \_152_[2] ;
 wire \_152_[30] ;
 wire \_152_[31] ;
 wire \_152_[3] ;
 wire \_152_[4] ;
 wire \_152_[5] ;
 wire \_152_[6] ;
 wire \_152_[7] ;
 wire \_152_[8] ;
 wire \_152_[9] ;
 wire \_158_[0] ;
 wire \_158_[10] ;
 wire \_158_[11] ;
 wire \_158_[12] ;
 wire \_158_[13] ;
 wire \_158_[14] ;
 wire \_158_[15] ;
 wire \_158_[16] ;
 wire \_158_[17] ;
 wire \_158_[18] ;
 wire \_158_[19] ;
 wire \_158_[1] ;
 wire \_158_[20] ;
 wire \_158_[21] ;
 wire \_158_[2] ;
 wire \_158_[3] ;
 wire \_158_[4] ;
 wire \_158_[5] ;
 wire \_158_[6] ;
 wire \_158_[7] ;
 wire \_158_[8] ;
 wire \_158_[9] ;
 wire \_164_[0] ;
 wire \_164_[10] ;
 wire \_164_[11] ;
 wire \_164_[12] ;
 wire \_164_[13] ;
 wire \_164_[14] ;
 wire \_164_[15] ;
 wire \_164_[16] ;
 wire \_164_[17] ;
 wire \_164_[18] ;
 wire \_164_[19] ;
 wire \_164_[1] ;
 wire \_164_[20] ;
 wire \_164_[21] ;
 wire \_164_[22] ;
 wire \_164_[23] ;
 wire \_164_[24] ;
 wire \_164_[25] ;
 wire \_164_[26] ;
 wire \_164_[27] ;
 wire \_164_[28] ;
 wire \_164_[29] ;
 wire \_164_[2] ;
 wire \_164_[30] ;
 wire \_164_[31] ;
 wire \_164_[3] ;
 wire \_164_[4] ;
 wire \_164_[5] ;
 wire \_164_[6] ;
 wire \_164_[7] ;
 wire \_164_[8] ;
 wire \_164_[9] ;
 wire \_167_[0] ;
 wire \_167_[10] ;
 wire \_167_[11] ;
 wire \_167_[12] ;
 wire \_167_[13] ;
 wire \_167_[14] ;
 wire \_167_[15] ;
 wire \_167_[16] ;
 wire \_167_[17] ;
 wire \_167_[18] ;
 wire \_167_[19] ;
 wire \_167_[1] ;
 wire \_167_[20] ;
 wire \_167_[21] ;
 wire \_167_[22] ;
 wire \_167_[23] ;
 wire \_167_[24] ;
 wire \_167_[25] ;
 wire \_167_[26] ;
 wire \_167_[27] ;
 wire \_167_[28] ;
 wire \_167_[29] ;
 wire \_167_[2] ;
 wire \_167_[30] ;
 wire \_167_[31] ;
 wire \_167_[3] ;
 wire \_167_[4] ;
 wire \_167_[5] ;
 wire \_167_[6] ;
 wire \_167_[7] ;
 wire \_167_[8] ;
 wire \_167_[9] ;
 wire \_170_[0] ;
 wire \_170_[10] ;
 wire \_170_[11] ;
 wire \_170_[12] ;
 wire \_170_[13] ;
 wire \_170_[14] ;
 wire \_170_[15] ;
 wire \_170_[16] ;
 wire \_170_[17] ;
 wire \_170_[18] ;
 wire \_170_[19] ;
 wire \_170_[1] ;
 wire \_170_[20] ;
 wire \_170_[21] ;
 wire \_170_[22] ;
 wire \_170_[23] ;
 wire \_170_[24] ;
 wire \_170_[25] ;
 wire \_170_[26] ;
 wire \_170_[27] ;
 wire \_170_[28] ;
 wire \_170_[29] ;
 wire \_170_[2] ;
 wire \_170_[30] ;
 wire \_170_[31] ;
 wire \_170_[3] ;
 wire \_170_[4] ;
 wire \_170_[5] ;
 wire \_170_[6] ;
 wire \_170_[7] ;
 wire \_170_[8] ;
 wire \_170_[9] ;
 wire \_173_[0] ;
 wire \_173_[10] ;
 wire \_173_[11] ;
 wire \_173_[12] ;
 wire \_173_[13] ;
 wire \_173_[14] ;
 wire \_173_[15] ;
 wire \_173_[16] ;
 wire \_173_[17] ;
 wire \_173_[18] ;
 wire \_173_[19] ;
 wire \_173_[1] ;
 wire \_173_[20] ;
 wire \_173_[21] ;
 wire \_173_[22] ;
 wire \_173_[23] ;
 wire \_173_[24] ;
 wire \_173_[25] ;
 wire \_173_[26] ;
 wire \_173_[27] ;
 wire \_173_[28] ;
 wire \_173_[29] ;
 wire \_173_[2] ;
 wire \_173_[30] ;
 wire \_173_[31] ;
 wire \_173_[3] ;
 wire \_173_[4] ;
 wire \_173_[5] ;
 wire \_173_[6] ;
 wire \_173_[7] ;
 wire \_173_[8] ;
 wire \_173_[9] ;
 wire \_176_[0] ;
 wire \_176_[10] ;
 wire \_176_[11] ;
 wire \_176_[12] ;
 wire \_176_[13] ;
 wire \_176_[14] ;
 wire \_176_[15] ;
 wire \_176_[16] ;
 wire \_176_[17] ;
 wire \_176_[18] ;
 wire \_176_[19] ;
 wire \_176_[1] ;
 wire \_176_[20] ;
 wire \_176_[21] ;
 wire \_176_[22] ;
 wire \_176_[23] ;
 wire \_176_[24] ;
 wire \_176_[25] ;
 wire \_176_[26] ;
 wire \_176_[27] ;
 wire \_176_[28] ;
 wire \_176_[29] ;
 wire \_176_[2] ;
 wire \_176_[30] ;
 wire \_176_[31] ;
 wire \_176_[3] ;
 wire \_176_[4] ;
 wire \_176_[5] ;
 wire \_176_[6] ;
 wire \_176_[7] ;
 wire \_176_[8] ;
 wire \_176_[9] ;
 wire \_179_[0] ;
 wire \_179_[10] ;
 wire \_179_[11] ;
 wire \_179_[12] ;
 wire \_179_[13] ;
 wire \_179_[14] ;
 wire \_179_[15] ;
 wire \_179_[16] ;
 wire \_179_[17] ;
 wire \_179_[18] ;
 wire \_179_[19] ;
 wire \_179_[1] ;
 wire \_179_[20] ;
 wire \_179_[21] ;
 wire \_179_[22] ;
 wire \_179_[23] ;
 wire \_179_[24] ;
 wire \_179_[25] ;
 wire \_179_[26] ;
 wire \_179_[27] ;
 wire \_179_[28] ;
 wire \_179_[29] ;
 wire \_179_[2] ;
 wire \_179_[30] ;
 wire \_179_[31] ;
 wire \_179_[3] ;
 wire \_179_[4] ;
 wire \_179_[5] ;
 wire \_179_[6] ;
 wire \_179_[7] ;
 wire \_179_[8] ;
 wire \_179_[9] ;
 wire \_182_[0] ;
 wire \_182_[10] ;
 wire \_182_[11] ;
 wire \_182_[12] ;
 wire \_182_[13] ;
 wire \_182_[14] ;
 wire \_182_[15] ;
 wire \_182_[16] ;
 wire \_182_[17] ;
 wire \_182_[18] ;
 wire \_182_[19] ;
 wire \_182_[1] ;
 wire \_182_[20] ;
 wire \_182_[21] ;
 wire \_182_[22] ;
 wire \_182_[23] ;
 wire \_182_[24] ;
 wire \_182_[25] ;
 wire \_182_[26] ;
 wire \_182_[27] ;
 wire \_182_[28] ;
 wire \_182_[29] ;
 wire \_182_[2] ;
 wire \_182_[30] ;
 wire \_182_[31] ;
 wire \_182_[3] ;
 wire \_182_[4] ;
 wire \_182_[5] ;
 wire \_182_[6] ;
 wire \_182_[7] ;
 wire \_182_[8] ;
 wire \_182_[9] ;
 wire \_185_[0] ;
 wire \_185_[10] ;
 wire \_185_[11] ;
 wire \_185_[12] ;
 wire \_185_[13] ;
 wire \_185_[14] ;
 wire \_185_[15] ;
 wire \_185_[16] ;
 wire \_185_[17] ;
 wire \_185_[18] ;
 wire \_185_[19] ;
 wire \_185_[1] ;
 wire \_185_[20] ;
 wire \_185_[21] ;
 wire \_185_[22] ;
 wire \_185_[23] ;
 wire \_185_[24] ;
 wire \_185_[25] ;
 wire \_185_[26] ;
 wire \_185_[27] ;
 wire \_185_[28] ;
 wire \_185_[29] ;
 wire \_185_[2] ;
 wire \_185_[30] ;
 wire \_185_[31] ;
 wire \_185_[3] ;
 wire \_185_[4] ;
 wire \_185_[5] ;
 wire \_185_[6] ;
 wire \_185_[7] ;
 wire \_185_[8] ;
 wire \_185_[9] ;
 wire \_190_[0] ;
 wire \_190_[1] ;
 wire \_190_[2] ;
 wire \_190_[3] ;
 wire \_195_[0] ;
 wire \_195_[1] ;
 wire \_195_[2] ;
 wire \_195_[3] ;
 wire \_195_[4] ;
 wire \_195_[5] ;
 wire \_225_[0] ;
 wire \_225_[10] ;
 wire \_225_[11] ;
 wire \_225_[12] ;
 wire \_225_[13] ;
 wire \_225_[14] ;
 wire \_225_[15] ;
 wire \_225_[16] ;
 wire \_225_[17] ;
 wire \_225_[18] ;
 wire \_225_[19] ;
 wire \_225_[1] ;
 wire \_225_[20] ;
 wire \_225_[21] ;
 wire \_225_[22] ;
 wire \_225_[23] ;
 wire \_225_[24] ;
 wire \_225_[25] ;
 wire \_225_[26] ;
 wire \_225_[27] ;
 wire \_225_[28] ;
 wire \_225_[29] ;
 wire \_225_[2] ;
 wire \_225_[30] ;
 wire \_225_[31] ;
 wire \_225_[3] ;
 wire \_225_[4] ;
 wire \_225_[5] ;
 wire \_225_[6] ;
 wire \_225_[7] ;
 wire \_225_[8] ;
 wire \_225_[9] ;
 wire \_228_[0] ;
 wire \_228_[10] ;
 wire \_228_[11] ;
 wire \_228_[12] ;
 wire \_228_[13] ;
 wire \_228_[14] ;
 wire \_228_[15] ;
 wire \_228_[16] ;
 wire \_228_[17] ;
 wire \_228_[18] ;
 wire \_228_[19] ;
 wire \_228_[1] ;
 wire \_228_[20] ;
 wire \_228_[21] ;
 wire \_228_[22] ;
 wire \_228_[23] ;
 wire \_228_[24] ;
 wire \_228_[25] ;
 wire \_228_[26] ;
 wire \_228_[27] ;
 wire \_228_[28] ;
 wire \_228_[29] ;
 wire \_228_[2] ;
 wire \_228_[30] ;
 wire \_228_[31] ;
 wire \_228_[3] ;
 wire \_228_[4] ;
 wire \_228_[5] ;
 wire \_228_[6] ;
 wire \_228_[7] ;
 wire \_228_[8] ;
 wire \_228_[9] ;
 wire \_231_[0] ;
 wire \_231_[10] ;
 wire \_231_[11] ;
 wire \_231_[12] ;
 wire \_231_[13] ;
 wire \_231_[14] ;
 wire \_231_[15] ;
 wire \_231_[16] ;
 wire \_231_[17] ;
 wire \_231_[18] ;
 wire \_231_[19] ;
 wire \_231_[1] ;
 wire \_231_[20] ;
 wire \_231_[21] ;
 wire \_231_[22] ;
 wire \_231_[23] ;
 wire \_231_[24] ;
 wire \_231_[25] ;
 wire \_231_[26] ;
 wire \_231_[27] ;
 wire \_231_[28] ;
 wire \_231_[29] ;
 wire \_231_[2] ;
 wire \_231_[30] ;
 wire \_231_[31] ;
 wire \_231_[3] ;
 wire \_231_[4] ;
 wire \_231_[5] ;
 wire \_231_[6] ;
 wire \_231_[7] ;
 wire \_231_[8] ;
 wire \_231_[9] ;
 wire \_234_[0] ;
 wire \_234_[10] ;
 wire \_234_[11] ;
 wire \_234_[12] ;
 wire \_234_[13] ;
 wire \_234_[14] ;
 wire \_234_[15] ;
 wire \_234_[16] ;
 wire \_234_[17] ;
 wire \_234_[18] ;
 wire \_234_[19] ;
 wire \_234_[1] ;
 wire \_234_[20] ;
 wire \_234_[21] ;
 wire \_234_[22] ;
 wire \_234_[23] ;
 wire \_234_[24] ;
 wire \_234_[25] ;
 wire \_234_[26] ;
 wire \_234_[27] ;
 wire \_234_[28] ;
 wire \_234_[29] ;
 wire \_234_[2] ;
 wire \_234_[30] ;
 wire \_234_[31] ;
 wire \_234_[3] ;
 wire \_234_[4] ;
 wire \_234_[5] ;
 wire \_234_[6] ;
 wire \_234_[7] ;
 wire \_234_[8] ;
 wire \_234_[9] ;
 wire \_237_[0] ;
 wire \_237_[10] ;
 wire \_237_[11] ;
 wire \_237_[12] ;
 wire \_237_[13] ;
 wire \_237_[14] ;
 wire \_237_[15] ;
 wire \_237_[16] ;
 wire \_237_[17] ;
 wire \_237_[18] ;
 wire \_237_[19] ;
 wire \_237_[1] ;
 wire \_237_[20] ;
 wire \_237_[21] ;
 wire \_237_[22] ;
 wire \_237_[23] ;
 wire \_237_[24] ;
 wire \_237_[25] ;
 wire \_237_[26] ;
 wire \_237_[27] ;
 wire \_237_[28] ;
 wire \_237_[29] ;
 wire \_237_[2] ;
 wire \_237_[30] ;
 wire \_237_[31] ;
 wire \_237_[3] ;
 wire \_237_[4] ;
 wire \_237_[5] ;
 wire \_237_[6] ;
 wire \_237_[7] ;
 wire \_237_[8] ;
 wire \_237_[9] ;
 wire \_240_[0] ;
 wire \_240_[10] ;
 wire \_240_[11] ;
 wire \_240_[12] ;
 wire \_240_[13] ;
 wire \_240_[14] ;
 wire \_240_[15] ;
 wire \_240_[16] ;
 wire \_240_[17] ;
 wire \_240_[18] ;
 wire \_240_[19] ;
 wire \_240_[1] ;
 wire \_240_[20] ;
 wire \_240_[21] ;
 wire \_240_[22] ;
 wire \_240_[23] ;
 wire \_240_[24] ;
 wire \_240_[25] ;
 wire \_240_[26] ;
 wire \_240_[27] ;
 wire \_240_[28] ;
 wire \_240_[29] ;
 wire \_240_[2] ;
 wire \_240_[30] ;
 wire \_240_[31] ;
 wire \_240_[3] ;
 wire \_240_[4] ;
 wire \_240_[5] ;
 wire \_240_[6] ;
 wire \_240_[7] ;
 wire \_240_[8] ;
 wire \_240_[9] ;
 wire \_243_[0] ;
 wire \_243_[10] ;
 wire \_243_[11] ;
 wire \_243_[12] ;
 wire \_243_[13] ;
 wire \_243_[14] ;
 wire \_243_[15] ;
 wire \_243_[16] ;
 wire \_243_[17] ;
 wire \_243_[18] ;
 wire \_243_[19] ;
 wire \_243_[1] ;
 wire \_243_[20] ;
 wire \_243_[21] ;
 wire \_243_[22] ;
 wire \_243_[23] ;
 wire \_243_[24] ;
 wire \_243_[25] ;
 wire \_243_[26] ;
 wire \_243_[27] ;
 wire \_243_[28] ;
 wire \_243_[29] ;
 wire \_243_[2] ;
 wire \_243_[30] ;
 wire \_243_[31] ;
 wire \_243_[3] ;
 wire \_243_[4] ;
 wire \_243_[5] ;
 wire \_243_[6] ;
 wire \_243_[7] ;
 wire \_243_[8] ;
 wire \_243_[9] ;
 wire \_246_[0] ;
 wire \_246_[10] ;
 wire \_246_[11] ;
 wire \_246_[12] ;
 wire \_246_[13] ;
 wire \_246_[14] ;
 wire \_246_[15] ;
 wire \_246_[16] ;
 wire \_246_[17] ;
 wire \_246_[18] ;
 wire \_246_[19] ;
 wire \_246_[1] ;
 wire \_246_[20] ;
 wire \_246_[21] ;
 wire \_246_[22] ;
 wire \_246_[23] ;
 wire \_246_[24] ;
 wire \_246_[25] ;
 wire \_246_[26] ;
 wire \_246_[27] ;
 wire \_246_[28] ;
 wire \_246_[29] ;
 wire \_246_[2] ;
 wire \_246_[30] ;
 wire \_246_[31] ;
 wire \_246_[3] ;
 wire \_246_[4] ;
 wire \_246_[5] ;
 wire \_246_[6] ;
 wire \_246_[7] ;
 wire \_246_[8] ;
 wire \_246_[9] ;
 wire \_392_[0] ;
 wire \_392_[1] ;
 wire \_392_[2] ;
 wire \_392_[3] ;
 wire \_392_[4] ;
 wire \_436_[0] ;
 wire \_436_[1] ;
 wire \_436_[2] ;
 wire \_436_[3] ;
 wire \_436_[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_1_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_opt_1_0_clk;

 sky130_fd_sc_hd__or2_2 _06492_ (.A(\_392_[1] ),
    .B(\_392_[0] ),
    .X(_01206_));
 sky130_fd_sc_hd__buf_2 _06493_ (.A(\_392_[2] ),
    .X(_01207_));
 sky130_fd_sc_hd__buf_2 _06494_ (.A(\_392_[3] ),
    .X(_01208_));
 sky130_fd_sc_hd__inv_2 _06495_ (.A(\_392_[4] ),
    .Y(_01209_));
 sky130_fd_sc_hd__or3_1 _06496_ (.A(_01207_),
    .B(_01208_),
    .C(_01209_),
    .X(_01210_));
 sky130_fd_sc_hd__or2_1 _06497_ (.A(_01206_),
    .B(_01210_),
    .X(_01211_));
 sky130_fd_sc_hd__or2_2 _06498_ (.A(net33),
    .B(_01211_),
    .X(_01212_));
 sky130_fd_sc_hd__inv_2 _06499_ (.A(_01212_),
    .Y(_01213_));
 sky130_fd_sc_hd__buf_4 _06500_ (.A(_01213_),
    .X(_01214_));
 sky130_fd_sc_hd__buf_6 _06501_ (.A(_01214_),
    .X(_01215_));
 sky130_fd_sc_hd__buf_6 _06502_ (.A(_01215_),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 _06503_ (.A(_01212_),
    .X(_01216_));
 sky130_fd_sc_hd__buf_4 _06504_ (.A(_01216_),
    .X(_01217_));
 sky130_fd_sc_hd__buf_6 _06505_ (.A(_01217_),
    .X(_01218_));
 sky130_fd_sc_hd__or4b_1 _06506_ (.A(\_190_[2] ),
    .B(\_190_[1] ),
    .C(\_190_[0] ),
    .D_N(\_190_[3] ),
    .X(_01219_));
 sky130_fd_sc_hd__and4_1 _06507_ (.A(\_190_[2] ),
    .B(\_190_[1] ),
    .C(\_190_[0] ),
    .D(_01213_),
    .X(_01220_));
 sky130_fd_sc_hd__xor2_1 _06508_ (.A(\_190_[3] ),
    .B(_01220_),
    .X(_01221_));
 sky130_fd_sc_hd__o21a_1 _06509_ (.A1(_01218_),
    .A2(_01219_),
    .B1(_01221_),
    .X(_00700_));
 sky130_fd_sc_hd__inv_2 _06510_ (.A(_01220_),
    .Y(_01222_));
 sky130_fd_sc_hd__a31o_1 _06511_ (.A1(\_190_[1] ),
    .A2(\_190_[0] ),
    .A3(_01215_),
    .B1(\_190_[2] ),
    .X(_01223_));
 sky130_fd_sc_hd__and2_1 _06512_ (.A(_01222_),
    .B(_01223_),
    .X(_01224_));
 sky130_fd_sc_hd__clkbuf_1 _06513_ (.A(_01224_),
    .X(_00699_));
 sky130_fd_sc_hd__clkbuf_4 _06514_ (.A(_01214_),
    .X(_01225_));
 sky130_fd_sc_hd__buf_6 _06515_ (.A(_01225_),
    .X(_01226_));
 sky130_fd_sc_hd__nand2_1 _06516_ (.A(\_190_[0] ),
    .B(_01226_),
    .Y(_01227_));
 sky130_fd_sc_hd__xnor2_1 _06517_ (.A(\_190_[1] ),
    .B(_01227_),
    .Y(_00698_));
 sky130_fd_sc_hd__or2_1 _06518_ (.A(\_190_[0] ),
    .B(_01215_),
    .X(_01228_));
 sky130_fd_sc_hd__and3_1 _06519_ (.A(_01227_),
    .B(_01219_),
    .C(_01228_),
    .X(_01229_));
 sky130_fd_sc_hd__clkbuf_1 _06520_ (.A(_01229_),
    .X(_00697_));
 sky130_fd_sc_hd__buf_2 _06521_ (.A(\_195_[5] ),
    .X(_01230_));
 sky130_fd_sc_hd__buf_2 _06522_ (.A(_01230_),
    .X(_01231_));
 sky130_fd_sc_hd__buf_2 _06523_ (.A(_01231_),
    .X(_01232_));
 sky130_fd_sc_hd__clkbuf_4 _06524_ (.A(_01232_),
    .X(_01233_));
 sky130_fd_sc_hd__buf_2 _06525_ (.A(\_195_[4] ),
    .X(_01234_));
 sky130_fd_sc_hd__buf_2 _06526_ (.A(_01234_),
    .X(_01235_));
 sky130_fd_sc_hd__buf_2 _06527_ (.A(_01235_),
    .X(_01236_));
 sky130_fd_sc_hd__buf_2 _06528_ (.A(_01236_),
    .X(_01237_));
 sky130_fd_sc_hd__buf_2 _06529_ (.A(_01237_),
    .X(_01238_));
 sky130_fd_sc_hd__clkbuf_4 _06530_ (.A(_01238_),
    .X(_01239_));
 sky130_fd_sc_hd__buf_2 _06531_ (.A(\_195_[3] ),
    .X(_01240_));
 sky130_fd_sc_hd__clkbuf_4 _06532_ (.A(_01240_),
    .X(_01241_));
 sky130_fd_sc_hd__buf_2 _06533_ (.A(_01241_),
    .X(_01242_));
 sky130_fd_sc_hd__buf_2 _06534_ (.A(_01242_),
    .X(_01243_));
 sky130_fd_sc_hd__buf_2 _06535_ (.A(_01243_),
    .X(_01244_));
 sky130_fd_sc_hd__or2b_1 _06536_ (.A(\_392_[3] ),
    .B_N(\_392_[2] ),
    .X(_01245_));
 sky130_fd_sc_hd__buf_2 _06537_ (.A(_01245_),
    .X(_01246_));
 sky130_fd_sc_hd__or3b_4 _06538_ (.A(_01207_),
    .B(\_392_[4] ),
    .C_N(_01208_),
    .X(_01247_));
 sky130_fd_sc_hd__or2_2 _06539_ (.A(_01206_),
    .B(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__o21ai_1 _06540_ (.A1(\_392_[4] ),
    .A2(_01246_),
    .B1(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__nand3_2 _06541_ (.A(\_392_[1] ),
    .B(\_392_[0] ),
    .C(_01209_),
    .Y(_01250_));
 sky130_fd_sc_hd__nand2_4 _06542_ (.A(_01207_),
    .B(_01208_),
    .Y(_01251_));
 sky130_fd_sc_hd__nor2_2 _06543_ (.A(_01250_),
    .B(_01251_),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_2 _06544_ (.A(_01249_),
    .B(_01252_),
    .Y(_01253_));
 sky130_fd_sc_hd__or4_2 _06545_ (.A(\_158_[1] ),
    .B(\_158_[0] ),
    .C(\_158_[3] ),
    .D(\_158_[2] ),
    .X(_01254_));
 sky130_fd_sc_hd__or3_1 _06546_ (.A(\_158_[5] ),
    .B(\_158_[4] ),
    .C(_01254_),
    .X(_01255_));
 sky130_fd_sc_hd__or2_2 _06547_ (.A(\_158_[6] ),
    .B(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__or3_1 _06548_ (.A(\_158_[7] ),
    .B(\_158_[8] ),
    .C(_01256_),
    .X(_01257_));
 sky130_fd_sc_hd__or2_1 _06549_ (.A(\_158_[9] ),
    .B(_01257_),
    .X(_01258_));
 sky130_fd_sc_hd__or3_1 _06550_ (.A(\_158_[11] ),
    .B(\_158_[10] ),
    .C(_01258_),
    .X(_01259_));
 sky130_fd_sc_hd__or2_1 _06551_ (.A(\_158_[12] ),
    .B(_01259_),
    .X(_01260_));
 sky130_fd_sc_hd__or3_1 _06552_ (.A(\_158_[13] ),
    .B(\_158_[14] ),
    .C(_01260_),
    .X(_01261_));
 sky130_fd_sc_hd__or2_1 _06553_ (.A(\_158_[15] ),
    .B(_01261_),
    .X(_01262_));
 sky130_fd_sc_hd__or3_1 _06554_ (.A(\_158_[17] ),
    .B(\_158_[16] ),
    .C(_01262_),
    .X(_01263_));
 sky130_fd_sc_hd__or2_1 _06555_ (.A(\_158_[18] ),
    .B(_01263_),
    .X(_01264_));
 sky130_fd_sc_hd__or3_1 _06556_ (.A(\_158_[19] ),
    .B(\_158_[20] ),
    .C(_01264_),
    .X(_01265_));
 sky130_fd_sc_hd__or2_2 _06557_ (.A(\_158_[21] ),
    .B(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__or3b_1 _06558_ (.A(\_392_[0] ),
    .B(\_392_[4] ),
    .C_N(\_392_[1] ),
    .X(_01267_));
 sky130_fd_sc_hd__buf_4 _06559_ (.A(_01267_),
    .X(_01268_));
 sky130_fd_sc_hd__nor2_8 _06560_ (.A(_01268_),
    .B(_01251_),
    .Y(_01269_));
 sky130_fd_sc_hd__or2_1 _06561_ (.A(_01252_),
    .B(_01269_),
    .X(_01270_));
 sky130_fd_sc_hd__a21oi_2 _06562_ (.A1(_01266_),
    .A2(_01270_),
    .B1(_01249_),
    .Y(_01271_));
 sky130_fd_sc_hd__or3_4 _06563_ (.A(\_392_[4] ),
    .B(_01206_),
    .C(_01251_),
    .X(_01272_));
 sky130_fd_sc_hd__nor2_1 _06564_ (.A(\_392_[1] ),
    .B(\_392_[0] ),
    .Y(_01273_));
 sky130_fd_sc_hd__or2_4 _06565_ (.A(_01273_),
    .B(_01247_),
    .X(_01274_));
 sky130_fd_sc_hd__o211a_1 _06566_ (.A1(net35),
    .A2(_01271_),
    .B1(_01272_),
    .C1(_01274_),
    .X(_01275_));
 sky130_fd_sc_hd__o21ai_4 _06567_ (.A1(net35),
    .A2(_01253_),
    .B1(_01275_),
    .Y(_01276_));
 sky130_fd_sc_hd__buf_2 _06568_ (.A(\_195_[2] ),
    .X(_01277_));
 sky130_fd_sc_hd__clkbuf_4 _06569_ (.A(_01277_),
    .X(_01278_));
 sky130_fd_sc_hd__buf_2 _06570_ (.A(\_195_[1] ),
    .X(_01279_));
 sky130_fd_sc_hd__clkbuf_4 _06571_ (.A(_01279_),
    .X(_01280_));
 sky130_fd_sc_hd__clkbuf_4 _06572_ (.A(_01280_),
    .X(_01281_));
 sky130_fd_sc_hd__clkbuf_4 _06573_ (.A(\_195_[0] ),
    .X(_01282_));
 sky130_fd_sc_hd__clkbuf_4 _06574_ (.A(_01282_),
    .X(_01283_));
 sky130_fd_sc_hd__clkbuf_4 _06575_ (.A(_01283_),
    .X(_01284_));
 sky130_fd_sc_hd__and3_1 _06576_ (.A(_01278_),
    .B(_01281_),
    .C(_01284_),
    .X(_01285_));
 sky130_fd_sc_hd__and3_1 _06577_ (.A(_01244_),
    .B(_01276_),
    .C(_01285_),
    .X(_01286_));
 sky130_fd_sc_hd__nand2_1 _06578_ (.A(_01239_),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__xnor2_1 _06579_ (.A(_01233_),
    .B(_01287_),
    .Y(_00408_));
 sky130_fd_sc_hd__or2_1 _06580_ (.A(_01239_),
    .B(_01286_),
    .X(_01288_));
 sky130_fd_sc_hd__and2_1 _06581_ (.A(_01287_),
    .B(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__clkbuf_1 _06582_ (.A(_01289_),
    .X(_00407_));
 sky130_fd_sc_hd__a21oi_1 _06583_ (.A1(_01276_),
    .A2(_01285_),
    .B1(_01244_),
    .Y(_01290_));
 sky130_fd_sc_hd__nor2_1 _06584_ (.A(_01286_),
    .B(_01290_),
    .Y(_00406_));
 sky130_fd_sc_hd__and2_1 _06585_ (.A(\_195_[1] ),
    .B(\_195_[0] ),
    .X(_01291_));
 sky130_fd_sc_hd__clkbuf_4 _06586_ (.A(_01291_),
    .X(_01292_));
 sky130_fd_sc_hd__a21oi_1 _06587_ (.A1(_01276_),
    .A2(_01292_),
    .B1(_01278_),
    .Y(_01293_));
 sky130_fd_sc_hd__a21oi_1 _06588_ (.A1(_01276_),
    .A2(_01285_),
    .B1(_01293_),
    .Y(_00405_));
 sky130_fd_sc_hd__a21oi_1 _06589_ (.A1(_01284_),
    .A2(_01276_),
    .B1(_01281_),
    .Y(_01294_));
 sky130_fd_sc_hd__a21oi_1 _06590_ (.A1(_01276_),
    .A2(_01292_),
    .B1(_01294_),
    .Y(_00404_));
 sky130_fd_sc_hd__clkbuf_4 _06591_ (.A(net35),
    .X(_01295_));
 sky130_fd_sc_hd__o21a_1 _06592_ (.A1(_01295_),
    .A2(_01253_),
    .B1(_01275_),
    .X(_01296_));
 sky130_fd_sc_hd__xnor2_1 _06593_ (.A(_01284_),
    .B(_01296_),
    .Y(_00403_));
 sky130_fd_sc_hd__nor2_2 _06594_ (.A(\_158_[21] ),
    .B(_01265_),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_1 _06595_ (.A(_099_),
    .B(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__or2_2 _06596_ (.A(_01268_),
    .B(_01251_),
    .X(_01299_));
 sky130_fd_sc_hd__clkbuf_2 _06597_ (.A(_01299_),
    .X(_01300_));
 sky130_fd_sc_hd__clkbuf_2 _06598_ (.A(_01300_),
    .X(_01301_));
 sky130_fd_sc_hd__buf_4 _06599_ (.A(_01301_),
    .X(_01302_));
 sky130_fd_sc_hd__inv_2 _06600_ (.A(net35),
    .Y(_01303_));
 sky130_fd_sc_hd__nor2_1 _06601_ (.A(_01303_),
    .B(_01297_),
    .Y(_01304_));
 sky130_fd_sc_hd__nor2_1 _06602_ (.A(_01302_),
    .B(_01304_),
    .Y(_01305_));
 sky130_fd_sc_hd__or3b_2 _06603_ (.A(\_392_[1] ),
    .B(\_392_[4] ),
    .C_N(\_392_[0] ),
    .X(_01306_));
 sky130_fd_sc_hd__or2_2 _06604_ (.A(_01306_),
    .B(_01251_),
    .X(_01307_));
 sky130_fd_sc_hd__nor2_1 _06605_ (.A(_01297_),
    .B(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__inv_2 _06606_ (.A(_01308_),
    .Y(_01309_));
 sky130_fd_sc_hd__or2_1 _06607_ (.A(_01208_),
    .B(_01306_),
    .X(_01310_));
 sky130_fd_sc_hd__o211a_1 _06608_ (.A1(_01208_),
    .A2(_01250_),
    .B1(_01310_),
    .C1(_01295_),
    .X(_01311_));
 sky130_fd_sc_hd__nor2_1 _06609_ (.A(_01246_),
    .B(_01268_),
    .Y(_01312_));
 sky130_fd_sc_hd__or3_4 _06610_ (.A(\_392_[4] ),
    .B(_01206_),
    .C(_01246_),
    .X(_01313_));
 sky130_fd_sc_hd__buf_2 _06611_ (.A(_01313_),
    .X(_01314_));
 sky130_fd_sc_hd__buf_2 _06612_ (.A(_01314_),
    .X(_01315_));
 sky130_fd_sc_hd__clkbuf_4 _06613_ (.A(_01315_),
    .X(_01316_));
 sky130_fd_sc_hd__inv_2 _06614_ (.A(_01316_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2_2 _06615_ (.A(_01206_),
    .B(_01247_),
    .Y(_01318_));
 sky130_fd_sc_hd__a211o_1 _06616_ (.A1(_093_),
    .A2(_01312_),
    .B1(_01317_),
    .C1(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__o2bb2a_1 _06617_ (.A1_N(_01309_),
    .A2_N(_01311_),
    .B1(_01319_),
    .B2(_01295_),
    .X(_01320_));
 sky130_fd_sc_hd__and3b_1 _06618_ (.A_N(_01251_),
    .B(_01209_),
    .C(_01273_),
    .X(_01321_));
 sky130_fd_sc_hd__a31o_1 _06619_ (.A1(\_392_[1] ),
    .A2(_01207_),
    .A3(_01209_),
    .B1(_01318_),
    .X(_01322_));
 sky130_fd_sc_hd__o21ba_1 _06620_ (.A1(_01246_),
    .A2(_01306_),
    .B1_N(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__or3_2 _06621_ (.A(_01207_),
    .B(_01208_),
    .C(_01250_),
    .X(_01324_));
 sky130_fd_sc_hd__or2_2 _06622_ (.A(_01207_),
    .B(_01310_),
    .X(_01325_));
 sky130_fd_sc_hd__nand3_1 _06623_ (.A(_01247_),
    .B(_01272_),
    .C(_01307_),
    .Y(_01326_));
 sky130_fd_sc_hd__o21ai_1 _06624_ (.A1(_01246_),
    .A2(_01306_),
    .B1(_01316_),
    .Y(_01327_));
 sky130_fd_sc_hd__nor3_1 _06625_ (.A(_01207_),
    .B(_01208_),
    .C(_01268_),
    .Y(_01328_));
 sky130_fd_sc_hd__a21oi_1 _06626_ (.A1(\_392_[1] ),
    .A2(\_392_[0] ),
    .B1(_01210_),
    .Y(_01329_));
 sky130_fd_sc_hd__or4_1 _06627_ (.A(net35),
    .B(_01327_),
    .C(_01328_),
    .D(_01329_),
    .X(_01330_));
 sky130_fd_sc_hd__nor2_1 _06628_ (.A(_01326_),
    .B(_01330_),
    .Y(_01331_));
 sky130_fd_sc_hd__and4_1 _06629_ (.A(_01323_),
    .B(_01324_),
    .C(_01325_),
    .D(_01331_),
    .X(_01332_));
 sky130_fd_sc_hd__nand2_1 _06630_ (.A(_099_),
    .B(_01295_),
    .Y(_01333_));
 sky130_fd_sc_hd__o21ai_1 _06631_ (.A1(_096_),
    .A2(_01306_),
    .B1(_01268_),
    .Y(_01334_));
 sky130_fd_sc_hd__and3b_1 _06632_ (.A_N(_01207_),
    .B(_01208_),
    .C(_01334_),
    .X(_01335_));
 sky130_fd_sc_hd__a221o_1 _06633_ (.A1(_01206_),
    .A2(_01329_),
    .B1(_01333_),
    .B2(_01328_),
    .C1(_01335_),
    .X(_01336_));
 sky130_fd_sc_hd__a2111o_1 _06634_ (.A1(_01295_),
    .A2(_01252_),
    .B1(_01321_),
    .C1(_01332_),
    .D1(_01336_),
    .X(_01337_));
 sky130_fd_sc_hd__a211o_1 _06635_ (.A1(_01298_),
    .A2(_01305_),
    .B1(_01320_),
    .C1(_01337_),
    .X(\_436_[0] ));
 sky130_fd_sc_hd__nor2_1 _06636_ (.A(_01304_),
    .B(_01307_),
    .Y(_01338_));
 sky130_fd_sc_hd__buf_4 _06637_ (.A(_01302_),
    .X(_01339_));
 sky130_fd_sc_hd__nor2_1 _06638_ (.A(_01297_),
    .B(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__or2_1 _06639_ (.A(_01252_),
    .B(_01340_),
    .X(_01341_));
 sky130_fd_sc_hd__nor2_1 _06640_ (.A(_01246_),
    .B(_01250_),
    .Y(_01342_));
 sky130_fd_sc_hd__a21o_1 _06641_ (.A1(_01295_),
    .A2(_01342_),
    .B1(_01312_),
    .X(_01343_));
 sky130_fd_sc_hd__nand2_1 _06642_ (.A(_096_),
    .B(_01208_),
    .Y(_01344_));
 sky130_fd_sc_hd__o21a_1 _06643_ (.A1(_01306_),
    .A2(_01344_),
    .B1(_01268_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _06644_ (.A0(_01310_),
    .A1(_01324_),
    .S(_01295_),
    .X(_01346_));
 sky130_fd_sc_hd__o221a_1 _06645_ (.A1(\_190_[3] ),
    .A2(_01222_),
    .B1(_01345_),
    .B2(_01207_),
    .C1(_01346_),
    .X(_01347_));
 sky130_fd_sc_hd__or4b_1 _06646_ (.A(_01338_),
    .B(_01341_),
    .C(_01343_),
    .D_N(_01347_),
    .X(_01348_));
 sky130_fd_sc_hd__clkbuf_1 _06647_ (.A(_01348_),
    .X(\_436_[1] ));
 sky130_fd_sc_hd__or3b_1 _06648_ (.A(_01250_),
    .B(_01207_),
    .C_N(_01208_),
    .X(_01349_));
 sky130_fd_sc_hd__o2111a_1 _06649_ (.A1(_01295_),
    .A2(_01324_),
    .B1(_01349_),
    .C1(_01272_),
    .D1(_01307_),
    .X(_01350_));
 sky130_fd_sc_hd__or4b_1 _06650_ (.A(_01327_),
    .B(_01343_),
    .C(_01341_),
    .D_N(_01350_),
    .X(_01351_));
 sky130_fd_sc_hd__clkbuf_1 _06651_ (.A(_01351_),
    .X(\_436_[2] ));
 sky130_fd_sc_hd__a21o_1 _06652_ (.A1(_01295_),
    .A2(_01252_),
    .B1(_01326_),
    .X(_01352_));
 sky130_fd_sc_hd__a211o_1 _06653_ (.A1(_01303_),
    .A2(_01342_),
    .B1(_01340_),
    .C1(_01352_),
    .X(\_436_[3] ));
 sky130_fd_sc_hd__buf_4 _06654_ (.A(_01302_),
    .X(_01353_));
 sky130_fd_sc_hd__buf_6 _06655_ (.A(_01353_),
    .X(_01354_));
 sky130_fd_sc_hd__buf_6 _06656_ (.A(_01354_),
    .X(_01355_));
 sky130_fd_sc_hd__o21ai_1 _06657_ (.A1(_01266_),
    .A2(_01355_),
    .B1(_01211_),
    .Y(\_436_[4] ));
 sky130_fd_sc_hd__nand2_1 _06658_ (.A(_099_),
    .B(_01328_),
    .Y(_01356_));
 sky130_fd_sc_hd__nand4_1 _06659_ (.A(_01253_),
    .B(_01324_),
    .C(_01325_),
    .D(_01356_),
    .Y(_01357_));
 sky130_fd_sc_hd__o31a_1 _06660_ (.A1(_01308_),
    .A2(_01340_),
    .A3(_01357_),
    .B1(_01303_),
    .X(net69));
 sky130_fd_sc_hd__nor2_4 _06661_ (.A(_01273_),
    .B(_01247_),
    .Y(_01358_));
 sky130_fd_sc_hd__a41o_1 _06662_ (.A1(_01302_),
    .A2(_01253_),
    .A3(_01309_),
    .A4(_01324_),
    .B1(net35),
    .X(_01359_));
 sky130_fd_sc_hd__or3b_2 _06663_ (.A(_01321_),
    .B(_01358_),
    .C_N(_01359_),
    .X(_01360_));
 sky130_fd_sc_hd__buf_4 _06664_ (.A(_01360_),
    .X(_01361_));
 sky130_fd_sc_hd__buf_4 _06665_ (.A(_01361_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _06666_ (.A0(\_116_[0] ),
    .A1(\_118_[0] ),
    .S(_01362_),
    .X(_01363_));
 sky130_fd_sc_hd__clkbuf_1 _06667_ (.A(_01363_),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _06668_ (.A0(\_116_[1] ),
    .A1(\_118_[1] ),
    .S(_01362_),
    .X(_01364_));
 sky130_fd_sc_hd__clkbuf_1 _06669_ (.A(_01364_),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _06670_ (.A0(\_116_[2] ),
    .A1(\_118_[2] ),
    .S(_01362_),
    .X(_01365_));
 sky130_fd_sc_hd__clkbuf_1 _06671_ (.A(_01365_),
    .X(_00117_));
 sky130_fd_sc_hd__and3_2 _06672_ (.A(_01272_),
    .B(_01274_),
    .C(_01359_),
    .X(_01366_));
 sky130_fd_sc_hd__buf_4 _06673_ (.A(_01366_),
    .X(_01367_));
 sky130_fd_sc_hd__buf_4 _06674_ (.A(_01367_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _06675_ (.A0(\_118_[3] ),
    .A1(\_116_[3] ),
    .S(_01368_),
    .X(_01369_));
 sky130_fd_sc_hd__clkbuf_1 _06676_ (.A(_01369_),
    .X(_00118_));
 sky130_fd_sc_hd__buf_4 _06677_ (.A(_01367_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _06678_ (.A0(\_118_[4] ),
    .A1(\_116_[4] ),
    .S(_01370_),
    .X(_01371_));
 sky130_fd_sc_hd__clkbuf_1 _06679_ (.A(_01371_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _06680_ (.A0(\_118_[5] ),
    .A1(\_116_[5] ),
    .S(_01370_),
    .X(_01372_));
 sky130_fd_sc_hd__clkbuf_1 _06681_ (.A(_01372_),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _06682_ (.A0(\_118_[6] ),
    .A1(\_116_[6] ),
    .S(_01370_),
    .X(_01373_));
 sky130_fd_sc_hd__clkbuf_1 _06683_ (.A(_01373_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _06684_ (.A0(\_118_[7] ),
    .A1(\_116_[7] ),
    .S(_01370_),
    .X(_01374_));
 sky130_fd_sc_hd__clkbuf_1 _06685_ (.A(_01374_),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _06686_ (.A0(\_118_[8] ),
    .A1(\_116_[8] ),
    .S(_01370_),
    .X(_01375_));
 sky130_fd_sc_hd__clkbuf_1 _06687_ (.A(_01375_),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _06688_ (.A0(\_118_[9] ),
    .A1(\_116_[9] ),
    .S(_01370_),
    .X(_01376_));
 sky130_fd_sc_hd__clkbuf_1 _06689_ (.A(_01376_),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _06690_ (.A0(\_118_[10] ),
    .A1(\_116_[10] ),
    .S(_01370_),
    .X(_01377_));
 sky130_fd_sc_hd__clkbuf_1 _06691_ (.A(_01377_),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _06692_ (.A0(\_118_[11] ),
    .A1(\_116_[11] ),
    .S(_01370_),
    .X(_01378_));
 sky130_fd_sc_hd__clkbuf_1 _06693_ (.A(_01378_),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _06694_ (.A0(\_118_[12] ),
    .A1(\_116_[12] ),
    .S(_01370_),
    .X(_01379_));
 sky130_fd_sc_hd__clkbuf_1 _06695_ (.A(_01379_),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _06696_ (.A0(\_118_[13] ),
    .A1(\_116_[13] ),
    .S(_01370_),
    .X(_01380_));
 sky130_fd_sc_hd__clkbuf_1 _06697_ (.A(_01380_),
    .X(_00128_));
 sky130_fd_sc_hd__buf_4 _06698_ (.A(_01367_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _06699_ (.A0(\_118_[14] ),
    .A1(\_116_[14] ),
    .S(_01381_),
    .X(_01382_));
 sky130_fd_sc_hd__clkbuf_1 _06700_ (.A(_01382_),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _06701_ (.A0(\_118_[15] ),
    .A1(\_116_[15] ),
    .S(_01381_),
    .X(_01383_));
 sky130_fd_sc_hd__clkbuf_1 _06702_ (.A(_01383_),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _06703_ (.A0(\_118_[16] ),
    .A1(\_116_[16] ),
    .S(_01381_),
    .X(_01384_));
 sky130_fd_sc_hd__clkbuf_1 _06704_ (.A(_01384_),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _06705_ (.A0(\_118_[17] ),
    .A1(\_116_[17] ),
    .S(_01381_),
    .X(_01385_));
 sky130_fd_sc_hd__clkbuf_1 _06706_ (.A(_01385_),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _06707_ (.A0(\_118_[18] ),
    .A1(\_116_[18] ),
    .S(_01381_),
    .X(_01386_));
 sky130_fd_sc_hd__clkbuf_1 _06708_ (.A(_01386_),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _06709_ (.A0(\_118_[19] ),
    .A1(\_116_[19] ),
    .S(_01381_),
    .X(_01387_));
 sky130_fd_sc_hd__clkbuf_1 _06710_ (.A(_01387_),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _06711_ (.A0(\_118_[20] ),
    .A1(\_116_[20] ),
    .S(_01381_),
    .X(_01388_));
 sky130_fd_sc_hd__clkbuf_1 _06712_ (.A(_01388_),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _06713_ (.A0(\_118_[21] ),
    .A1(\_116_[21] ),
    .S(_01381_),
    .X(_01389_));
 sky130_fd_sc_hd__clkbuf_1 _06714_ (.A(_01389_),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _06715_ (.A0(\_118_[22] ),
    .A1(\_116_[22] ),
    .S(_01381_),
    .X(_01390_));
 sky130_fd_sc_hd__clkbuf_1 _06716_ (.A(_01390_),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _06717_ (.A0(\_118_[23] ),
    .A1(\_116_[23] ),
    .S(_01381_),
    .X(_01391_));
 sky130_fd_sc_hd__clkbuf_1 _06718_ (.A(_01391_),
    .X(_00138_));
 sky130_fd_sc_hd__buf_4 _06719_ (.A(_01366_),
    .X(_01392_));
 sky130_fd_sc_hd__clkbuf_4 _06720_ (.A(_01392_),
    .X(_01393_));
 sky130_fd_sc_hd__buf_4 _06721_ (.A(_01393_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _06722_ (.A0(\_118_[24] ),
    .A1(\_116_[24] ),
    .S(_01394_),
    .X(_01395_));
 sky130_fd_sc_hd__clkbuf_1 _06723_ (.A(_01395_),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _06724_ (.A0(\_118_[25] ),
    .A1(\_116_[25] ),
    .S(_01394_),
    .X(_01396_));
 sky130_fd_sc_hd__clkbuf_1 _06725_ (.A(_01396_),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _06726_ (.A0(\_118_[26] ),
    .A1(\_116_[26] ),
    .S(_01394_),
    .X(_01397_));
 sky130_fd_sc_hd__clkbuf_1 _06727_ (.A(_01397_),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _06728_ (.A0(\_118_[27] ),
    .A1(\_116_[27] ),
    .S(_01394_),
    .X(_01398_));
 sky130_fd_sc_hd__clkbuf_1 _06729_ (.A(_01398_),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _06730_ (.A0(\_118_[28] ),
    .A1(\_116_[28] ),
    .S(_01394_),
    .X(_01399_));
 sky130_fd_sc_hd__clkbuf_1 _06731_ (.A(_01399_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _06732_ (.A0(\_118_[29] ),
    .A1(\_116_[29] ),
    .S(_01394_),
    .X(_01400_));
 sky130_fd_sc_hd__clkbuf_1 _06733_ (.A(_01400_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _06734_ (.A0(\_118_[30] ),
    .A1(\_116_[30] ),
    .S(_01394_),
    .X(_01401_));
 sky130_fd_sc_hd__clkbuf_1 _06735_ (.A(_01401_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _06736_ (.A0(\_118_[31] ),
    .A1(\_116_[31] ),
    .S(_01394_),
    .X(_01402_));
 sky130_fd_sc_hd__clkbuf_1 _06737_ (.A(_01402_),
    .X(_00146_));
 sky130_fd_sc_hd__inv_2 _06738_ (.A(net34),
    .Y(_00100_));
 sky130_fd_sc_hd__inv_2 _06739_ (.A(net34),
    .Y(_00101_));
 sky130_fd_sc_hd__inv_2 _06740_ (.A(net34),
    .Y(_00102_));
 sky130_fd_sc_hd__inv_2 _06741_ (.A(net34),
    .Y(_00103_));
 sky130_fd_sc_hd__inv_2 _06742_ (.A(net34),
    .Y(_00104_));
 sky130_fd_sc_hd__a21oi_2 _06743_ (.A1(_01323_),
    .A2(_01307_),
    .B1(_01304_),
    .Y(_01403_));
 sky130_fd_sc_hd__nor3_4 _06744_ (.A(_01321_),
    .B(_01358_),
    .C(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__buf_4 _06745_ (.A(_01404_),
    .X(_01405_));
 sky130_fd_sc_hd__buf_4 _06746_ (.A(_01405_),
    .X(_01406_));
 sky130_fd_sc_hd__clkbuf_4 _06747_ (.A(_01406_),
    .X(_01407_));
 sky130_fd_sc_hd__buf_4 _06748_ (.A(_01269_),
    .X(_01408_));
 sky130_fd_sc_hd__buf_4 _06749_ (.A(_01408_),
    .X(_01409_));
 sky130_fd_sc_hd__or3_1 _06750_ (.A(_01321_),
    .B(_01358_),
    .C(_01403_),
    .X(_01410_));
 sky130_fd_sc_hd__buf_6 _06751_ (.A(_01410_),
    .X(_01411_));
 sky130_fd_sc_hd__clkbuf_4 _06752_ (.A(_01411_),
    .X(_01412_));
 sky130_fd_sc_hd__or2_1 _06753_ (.A(\_179_[0] ),
    .B(_01299_),
    .X(_01413_));
 sky130_fd_sc_hd__o211a_1 _06754_ (.A1(\_243_[0] ),
    .A2(_01409_),
    .B1(_01412_),
    .C1(_01413_),
    .X(_01414_));
 sky130_fd_sc_hd__nor2_1 _06755_ (.A(\_392_[0] ),
    .B(_01210_),
    .Y(_01415_));
 sky130_fd_sc_hd__a21o_2 _06756_ (.A1(\_392_[1] ),
    .A2(_01415_),
    .B1(net34),
    .X(_01416_));
 sky130_fd_sc_hd__buf_4 _06757_ (.A(_01416_),
    .X(_01417_));
 sky130_fd_sc_hd__clkbuf_4 _06758_ (.A(_01417_),
    .X(_01418_));
 sky130_fd_sc_hd__buf_4 _06759_ (.A(_01418_),
    .X(_01419_));
 sky130_fd_sc_hd__a211o_1 _06760_ (.A1(\_246_[0] ),
    .A2(_01407_),
    .B1(_01414_),
    .C1(_01419_),
    .X(_00147_));
 sky130_fd_sc_hd__clkbuf_4 _06761_ (.A(_01411_),
    .X(_01420_));
 sky130_fd_sc_hd__clkbuf_8 _06762_ (.A(_01420_),
    .X(_01421_));
 sky130_fd_sc_hd__buf_2 _06763_ (.A(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__inv_2 _06764_ (.A(_01416_),
    .Y(_01423_));
 sky130_fd_sc_hd__buf_4 _06765_ (.A(_01423_),
    .X(_01424_));
 sky130_fd_sc_hd__clkbuf_4 _06766_ (.A(_01424_),
    .X(_01425_));
 sky130_fd_sc_hd__clkbuf_8 _06767_ (.A(_01412_),
    .X(_01426_));
 sky130_fd_sc_hd__buf_4 _06768_ (.A(_01408_),
    .X(_01427_));
 sky130_fd_sc_hd__buf_4 _06769_ (.A(_01427_),
    .X(_01428_));
 sky130_fd_sc_hd__or3_1 _06770_ (.A(\_179_[1] ),
    .B(_01268_),
    .C(_01251_),
    .X(_01429_));
 sky130_fd_sc_hd__o21ai_1 _06771_ (.A1(\_243_[1] ),
    .A2(_01428_),
    .B1(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__nand2_1 _06772_ (.A(_01426_),
    .B(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hd__o211a_1 _06773_ (.A1(\_246_[1] ),
    .A2(_01422_),
    .B1(_01425_),
    .C1(_01431_),
    .X(_00148_));
 sky130_fd_sc_hd__or3_1 _06774_ (.A(\_179_[2] ),
    .B(_01268_),
    .C(_01251_),
    .X(_01432_));
 sky130_fd_sc_hd__o21ai_1 _06775_ (.A1(\_243_[2] ),
    .A2(_01428_),
    .B1(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_1 _06776_ (.A(_01426_),
    .B(_01433_),
    .Y(_01434_));
 sky130_fd_sc_hd__o211a_1 _06777_ (.A1(\_246_[2] ),
    .A2(_01422_),
    .B1(_01425_),
    .C1(_01434_),
    .X(_00149_));
 sky130_fd_sc_hd__buf_4 _06778_ (.A(_01416_),
    .X(_01435_));
 sky130_fd_sc_hd__buf_4 _06779_ (.A(_01435_),
    .X(_01436_));
 sky130_fd_sc_hd__buf_4 _06780_ (.A(_01408_),
    .X(_01437_));
 sky130_fd_sc_hd__clkbuf_4 _06781_ (.A(_01437_),
    .X(_01438_));
 sky130_fd_sc_hd__buf_4 _06782_ (.A(_01411_),
    .X(_01439_));
 sky130_fd_sc_hd__or2_1 _06783_ (.A(\_179_[3] ),
    .B(_01299_),
    .X(_01440_));
 sky130_fd_sc_hd__o211a_1 _06784_ (.A1(\_243_[3] ),
    .A2(_01438_),
    .B1(_01439_),
    .C1(_01440_),
    .X(_01441_));
 sky130_fd_sc_hd__a211o_1 _06785_ (.A1(\_246_[3] ),
    .A2(_01407_),
    .B1(_01436_),
    .C1(_01441_),
    .X(_00150_));
 sky130_fd_sc_hd__or2_1 _06786_ (.A(\_179_[4] ),
    .B(_01299_),
    .X(_01442_));
 sky130_fd_sc_hd__o211a_1 _06787_ (.A1(\_243_[4] ),
    .A2(_01438_),
    .B1(_01439_),
    .C1(_01442_),
    .X(_01443_));
 sky130_fd_sc_hd__a211o_1 _06788_ (.A1(\_246_[4] ),
    .A2(_01407_),
    .B1(_01436_),
    .C1(_01443_),
    .X(_00151_));
 sky130_fd_sc_hd__clkbuf_4 _06789_ (.A(_01412_),
    .X(_01444_));
 sky130_fd_sc_hd__or2_1 _06790_ (.A(\_179_[5] ),
    .B(_01299_),
    .X(_01445_));
 sky130_fd_sc_hd__o21ai_1 _06791_ (.A1(\_243_[5] ),
    .A2(_01428_),
    .B1(_01445_),
    .Y(_01446_));
 sky130_fd_sc_hd__nand2_1 _06792_ (.A(_01444_),
    .B(_01446_),
    .Y(_01447_));
 sky130_fd_sc_hd__o211a_1 _06793_ (.A1(\_246_[5] ),
    .A2(_01422_),
    .B1(_01425_),
    .C1(_01447_),
    .X(_00152_));
 sky130_fd_sc_hd__buf_2 _06794_ (.A(_01405_),
    .X(_01448_));
 sky130_fd_sc_hd__buf_4 _06795_ (.A(_01339_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _06796_ (.A0(\_179_[6] ),
    .A1(\_243_[6] ),
    .S(_01449_),
    .X(_01450_));
 sky130_fd_sc_hd__or2_1 _06797_ (.A(_01448_),
    .B(_01450_),
    .X(_01451_));
 sky130_fd_sc_hd__o211a_1 _06798_ (.A1(\_246_[6] ),
    .A2(_01422_),
    .B1(_01425_),
    .C1(_01451_),
    .X(_00153_));
 sky130_fd_sc_hd__or2_1 _06799_ (.A(\_179_[7] ),
    .B(_01300_),
    .X(_01452_));
 sky130_fd_sc_hd__o21ai_1 _06800_ (.A1(\_243_[7] ),
    .A2(_01428_),
    .B1(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand2_1 _06801_ (.A(_01444_),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__o211a_1 _06802_ (.A1(\_246_[7] ),
    .A2(_01422_),
    .B1(_01425_),
    .C1(_01454_),
    .X(_00154_));
 sky130_fd_sc_hd__or2_1 _06803_ (.A(\_179_[8] ),
    .B(_01299_),
    .X(_01455_));
 sky130_fd_sc_hd__o211a_1 _06804_ (.A1(\_243_[8] ),
    .A2(_01438_),
    .B1(_01439_),
    .C1(_01455_),
    .X(_01456_));
 sky130_fd_sc_hd__a211o_1 _06805_ (.A1(\_246_[8] ),
    .A2(_01407_),
    .B1(_01436_),
    .C1(_01456_),
    .X(_00155_));
 sky130_fd_sc_hd__or2_1 _06806_ (.A(\_179_[9] ),
    .B(_01300_),
    .X(_01457_));
 sky130_fd_sc_hd__o21ai_1 _06807_ (.A1(\_243_[9] ),
    .A2(_01428_),
    .B1(_01457_),
    .Y(_01458_));
 sky130_fd_sc_hd__nand2_1 _06808_ (.A(_01444_),
    .B(_01458_),
    .Y(_01459_));
 sky130_fd_sc_hd__o211a_1 _06809_ (.A1(\_246_[9] ),
    .A2(_01422_),
    .B1(_01425_),
    .C1(_01459_),
    .X(_00156_));
 sky130_fd_sc_hd__buf_2 _06810_ (.A(_01435_),
    .X(_01460_));
 sky130_fd_sc_hd__buf_2 _06811_ (.A(_01420_),
    .X(_01461_));
 sky130_fd_sc_hd__or2_1 _06812_ (.A(\_179_[10] ),
    .B(_01300_),
    .X(_01462_));
 sky130_fd_sc_hd__o211a_1 _06813_ (.A1(\_243_[10] ),
    .A2(_01438_),
    .B1(_01461_),
    .C1(_01462_),
    .X(_01463_));
 sky130_fd_sc_hd__a211o_1 _06814_ (.A1(\_246_[10] ),
    .A2(_01407_),
    .B1(_01460_),
    .C1(_01463_),
    .X(_00157_));
 sky130_fd_sc_hd__or2_1 _06815_ (.A(\_179_[11] ),
    .B(_01299_),
    .X(_01464_));
 sky130_fd_sc_hd__o211a_1 _06816_ (.A1(\_243_[11] ),
    .A2(_01438_),
    .B1(_01461_),
    .C1(_01464_),
    .X(_01465_));
 sky130_fd_sc_hd__a211o_1 _06817_ (.A1(\_246_[11] ),
    .A2(_01407_),
    .B1(_01460_),
    .C1(_01465_),
    .X(_00158_));
 sky130_fd_sc_hd__or2_1 _06818_ (.A(\_179_[12] ),
    .B(_01299_),
    .X(_01466_));
 sky130_fd_sc_hd__o21ai_1 _06819_ (.A1(\_243_[12] ),
    .A2(_01428_),
    .B1(_01466_),
    .Y(_01467_));
 sky130_fd_sc_hd__nand2_1 _06820_ (.A(_01444_),
    .B(_01467_),
    .Y(_01468_));
 sky130_fd_sc_hd__o211a_1 _06821_ (.A1(\_246_[12] ),
    .A2(_01422_),
    .B1(_01425_),
    .C1(_01468_),
    .X(_00159_));
 sky130_fd_sc_hd__or2_1 _06822_ (.A(\_179_[13] ),
    .B(_01300_),
    .X(_01469_));
 sky130_fd_sc_hd__o21ai_1 _06823_ (.A1(\_243_[13] ),
    .A2(_01428_),
    .B1(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hd__nand2_1 _06824_ (.A(_01444_),
    .B(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hd__o211a_1 _06825_ (.A1(\_246_[13] ),
    .A2(_01422_),
    .B1(_01425_),
    .C1(_01471_),
    .X(_00160_));
 sky130_fd_sc_hd__or2_1 _06826_ (.A(\_179_[14] ),
    .B(_01300_),
    .X(_01472_));
 sky130_fd_sc_hd__o211a_1 _06827_ (.A1(\_243_[14] ),
    .A2(_01438_),
    .B1(_01461_),
    .C1(_01472_),
    .X(_01473_));
 sky130_fd_sc_hd__a211o_1 _06828_ (.A1(\_246_[14] ),
    .A2(_01407_),
    .B1(_01460_),
    .C1(_01473_),
    .X(_00161_));
 sky130_fd_sc_hd__clkbuf_4 _06829_ (.A(_01427_),
    .X(_01474_));
 sky130_fd_sc_hd__or2_1 _06830_ (.A(\_179_[15] ),
    .B(_01300_),
    .X(_01475_));
 sky130_fd_sc_hd__o211a_1 _06831_ (.A1(\_243_[15] ),
    .A2(_01474_),
    .B1(_01461_),
    .C1(_01475_),
    .X(_01476_));
 sky130_fd_sc_hd__a211o_1 _06832_ (.A1(\_246_[15] ),
    .A2(_01407_),
    .B1(_01460_),
    .C1(_01476_),
    .X(_00162_));
 sky130_fd_sc_hd__or2_1 _06833_ (.A(\_179_[16] ),
    .B(_01301_),
    .X(_01477_));
 sky130_fd_sc_hd__o21ai_1 _06834_ (.A1(\_243_[16] ),
    .A2(_01438_),
    .B1(_01477_),
    .Y(_01478_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(_01444_),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__o211a_1 _06836_ (.A1(\_246_[16] ),
    .A2(_01422_),
    .B1(_01425_),
    .C1(_01479_),
    .X(_00163_));
 sky130_fd_sc_hd__buf_4 _06837_ (.A(_01423_),
    .X(_01480_));
 sky130_fd_sc_hd__buf_2 _06838_ (.A(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__or2_1 _06839_ (.A(\_179_[17] ),
    .B(_01300_),
    .X(_01482_));
 sky130_fd_sc_hd__o21ai_1 _06840_ (.A1(\_243_[17] ),
    .A2(_01438_),
    .B1(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hd__nand2_1 _06841_ (.A(_01444_),
    .B(_01483_),
    .Y(_01484_));
 sky130_fd_sc_hd__o211a_1 _06842_ (.A1(\_246_[17] ),
    .A2(_01422_),
    .B1(_01481_),
    .C1(_01484_),
    .X(_00164_));
 sky130_fd_sc_hd__clkbuf_4 _06843_ (.A(_01421_),
    .X(_01485_));
 sky130_fd_sc_hd__or2_1 _06844_ (.A(\_179_[18] ),
    .B(_01300_),
    .X(_01486_));
 sky130_fd_sc_hd__o21ai_1 _06845_ (.A1(\_243_[18] ),
    .A2(_01438_),
    .B1(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hd__nand2_1 _06846_ (.A(_01444_),
    .B(_01487_),
    .Y(_01488_));
 sky130_fd_sc_hd__o211a_1 _06847_ (.A1(\_246_[18] ),
    .A2(_01485_),
    .B1(_01481_),
    .C1(_01488_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _06848_ (.A0(\_179_[19] ),
    .A1(\_243_[19] ),
    .S(_01449_),
    .X(_01489_));
 sky130_fd_sc_hd__or2_1 _06849_ (.A(_01448_),
    .B(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__o211a_1 _06850_ (.A1(\_246_[19] ),
    .A2(_01485_),
    .B1(_01481_),
    .C1(_01490_),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _06851_ (.A0(\_179_[20] ),
    .A1(\_243_[20] ),
    .S(_01449_),
    .X(_01491_));
 sky130_fd_sc_hd__or2_1 _06852_ (.A(_01448_),
    .B(_01491_),
    .X(_01492_));
 sky130_fd_sc_hd__o211a_1 _06853_ (.A1(\_246_[20] ),
    .A2(_01485_),
    .B1(_01481_),
    .C1(_01492_),
    .X(_00167_));
 sky130_fd_sc_hd__or2_1 _06854_ (.A(\_179_[21] ),
    .B(_01301_),
    .X(_01493_));
 sky130_fd_sc_hd__o211a_1 _06855_ (.A1(\_243_[21] ),
    .A2(_01474_),
    .B1(_01461_),
    .C1(_01493_),
    .X(_01494_));
 sky130_fd_sc_hd__a211o_1 _06856_ (.A1(\_246_[21] ),
    .A2(_01407_),
    .B1(_01460_),
    .C1(_01494_),
    .X(_00168_));
 sky130_fd_sc_hd__buf_4 _06857_ (.A(_01405_),
    .X(_01495_));
 sky130_fd_sc_hd__clkbuf_4 _06858_ (.A(_01495_),
    .X(_01496_));
 sky130_fd_sc_hd__or2_1 _06859_ (.A(\_179_[22] ),
    .B(_01301_),
    .X(_01497_));
 sky130_fd_sc_hd__o211a_1 _06860_ (.A1(\_243_[22] ),
    .A2(_01474_),
    .B1(_01461_),
    .C1(_01497_),
    .X(_01498_));
 sky130_fd_sc_hd__a211o_1 _06861_ (.A1(\_246_[22] ),
    .A2(_01496_),
    .B1(_01460_),
    .C1(_01498_),
    .X(_00169_));
 sky130_fd_sc_hd__or2_1 _06862_ (.A(\_179_[23] ),
    .B(_01301_),
    .X(_01499_));
 sky130_fd_sc_hd__o211a_1 _06863_ (.A1(\_243_[23] ),
    .A2(_01474_),
    .B1(_01461_),
    .C1(_01499_),
    .X(_01500_));
 sky130_fd_sc_hd__a211o_1 _06864_ (.A1(\_246_[23] ),
    .A2(_01496_),
    .B1(_01460_),
    .C1(_01500_),
    .X(_00170_));
 sky130_fd_sc_hd__or2_1 _06865_ (.A(\_179_[24] ),
    .B(_01301_),
    .X(_01501_));
 sky130_fd_sc_hd__o211a_1 _06866_ (.A1(\_243_[24] ),
    .A2(_01474_),
    .B1(_01461_),
    .C1(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__a211o_1 _06867_ (.A1(\_246_[24] ),
    .A2(_01496_),
    .B1(_01460_),
    .C1(_01502_),
    .X(_00171_));
 sky130_fd_sc_hd__or2_1 _06868_ (.A(\_179_[25] ),
    .B(_01301_),
    .X(_01503_));
 sky130_fd_sc_hd__o211a_1 _06869_ (.A1(\_243_[25] ),
    .A2(_01474_),
    .B1(_01461_),
    .C1(_01503_),
    .X(_01504_));
 sky130_fd_sc_hd__a211o_1 _06870_ (.A1(\_246_[25] ),
    .A2(_01496_),
    .B1(_01460_),
    .C1(_01504_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _06871_ (.A0(\_179_[26] ),
    .A1(\_243_[26] ),
    .S(_01449_),
    .X(_01505_));
 sky130_fd_sc_hd__or2_1 _06872_ (.A(_01448_),
    .B(_01505_),
    .X(_01506_));
 sky130_fd_sc_hd__o211a_1 _06873_ (.A1(\_246_[26] ),
    .A2(_01485_),
    .B1(_01481_),
    .C1(_01506_),
    .X(_00173_));
 sky130_fd_sc_hd__or2_1 _06874_ (.A(\_179_[27] ),
    .B(_01301_),
    .X(_01507_));
 sky130_fd_sc_hd__o211a_1 _06875_ (.A1(\_243_[27] ),
    .A2(_01474_),
    .B1(_01461_),
    .C1(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__a211o_1 _06876_ (.A1(\_246_[27] ),
    .A2(_01496_),
    .B1(_01460_),
    .C1(_01508_),
    .X(_00174_));
 sky130_fd_sc_hd__clkbuf_4 _06877_ (.A(_01435_),
    .X(_01509_));
 sky130_fd_sc_hd__buf_2 _06878_ (.A(_01420_),
    .X(_01510_));
 sky130_fd_sc_hd__or2_1 _06879_ (.A(\_179_[28] ),
    .B(_01302_),
    .X(_01511_));
 sky130_fd_sc_hd__o211a_1 _06880_ (.A1(\_243_[28] ),
    .A2(_01474_),
    .B1(_01510_),
    .C1(_01511_),
    .X(_01512_));
 sky130_fd_sc_hd__a211o_1 _06881_ (.A1(\_246_[28] ),
    .A2(_01496_),
    .B1(_01509_),
    .C1(_01512_),
    .X(_00175_));
 sky130_fd_sc_hd__or2_1 _06882_ (.A(\_179_[29] ),
    .B(_01302_),
    .X(_01513_));
 sky130_fd_sc_hd__o21ai_1 _06883_ (.A1(\_243_[29] ),
    .A2(_01438_),
    .B1(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__nand2_1 _06884_ (.A(_01444_),
    .B(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__o211a_1 _06885_ (.A1(\_246_[29] ),
    .A2(_01485_),
    .B1(_01481_),
    .C1(_01515_),
    .X(_00176_));
 sky130_fd_sc_hd__or2_1 _06886_ (.A(\_179_[30] ),
    .B(_01302_),
    .X(_01516_));
 sky130_fd_sc_hd__o211a_1 _06887_ (.A1(\_243_[30] ),
    .A2(_01474_),
    .B1(_01510_),
    .C1(_01516_),
    .X(_01517_));
 sky130_fd_sc_hd__a211o_1 _06888_ (.A1(\_246_[30] ),
    .A2(_01496_),
    .B1(_01509_),
    .C1(_01517_),
    .X(_00177_));
 sky130_fd_sc_hd__buf_4 _06889_ (.A(_01302_),
    .X(_01518_));
 sky130_fd_sc_hd__buf_4 _06890_ (.A(_01518_),
    .X(_01519_));
 sky130_fd_sc_hd__buf_4 _06891_ (.A(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__and2_1 _06892_ (.A(\_179_[31] ),
    .B(_01269_),
    .X(_01521_));
 sky130_fd_sc_hd__a211o_1 _06893_ (.A1(\_243_[31] ),
    .A2(_01520_),
    .B1(_01495_),
    .C1(_01521_),
    .X(_01522_));
 sky130_fd_sc_hd__o211a_1 _06894_ (.A1(\_246_[31] ),
    .A2(_01485_),
    .B1(_01481_),
    .C1(_01522_),
    .X(_00178_));
 sky130_fd_sc_hd__clkbuf_8 _06895_ (.A(_01353_),
    .X(_01523_));
 sky130_fd_sc_hd__or2_1 _06896_ (.A(\_176_[0] ),
    .B(_01523_),
    .X(_01524_));
 sky130_fd_sc_hd__o211a_1 _06897_ (.A1(\_240_[0] ),
    .A2(_01474_),
    .B1(_01510_),
    .C1(_01524_),
    .X(_01525_));
 sky130_fd_sc_hd__a211o_1 _06898_ (.A1(\_243_[0] ),
    .A2(_01496_),
    .B1(_01509_),
    .C1(_01525_),
    .X(_00179_));
 sky130_fd_sc_hd__clkbuf_4 _06899_ (.A(_01427_),
    .X(_01526_));
 sky130_fd_sc_hd__or2_1 _06900_ (.A(\_176_[1] ),
    .B(_01523_),
    .X(_01527_));
 sky130_fd_sc_hd__o211a_1 _06901_ (.A1(\_240_[1] ),
    .A2(_01526_),
    .B1(_01510_),
    .C1(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__a211o_1 _06902_ (.A1(\_243_[1] ),
    .A2(_01496_),
    .B1(_01509_),
    .C1(_01528_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _06903_ (.A0(\_176_[2] ),
    .A1(\_240_[2] ),
    .S(_01449_),
    .X(_01529_));
 sky130_fd_sc_hd__or2_1 _06904_ (.A(_01448_),
    .B(_01529_),
    .X(_01530_));
 sky130_fd_sc_hd__o211a_1 _06905_ (.A1(\_243_[2] ),
    .A2(_01485_),
    .B1(_01481_),
    .C1(_01530_),
    .X(_00181_));
 sky130_fd_sc_hd__clkbuf_2 _06906_ (.A(_01339_),
    .X(_01531_));
 sky130_fd_sc_hd__or2_1 _06907_ (.A(\_176_[3] ),
    .B(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__o211a_1 _06908_ (.A1(\_240_[3] ),
    .A2(_01526_),
    .B1(_01510_),
    .C1(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__a211o_1 _06909_ (.A1(\_243_[3] ),
    .A2(_01496_),
    .B1(_01509_),
    .C1(_01533_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _06910_ (.A0(\_176_[4] ),
    .A1(\_240_[4] ),
    .S(_01449_),
    .X(_01534_));
 sky130_fd_sc_hd__or2_1 _06911_ (.A(_01448_),
    .B(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__o211a_1 _06912_ (.A1(\_243_[4] ),
    .A2(_01485_),
    .B1(_01481_),
    .C1(_01535_),
    .X(_00183_));
 sky130_fd_sc_hd__clkbuf_4 _06913_ (.A(_01495_),
    .X(_01536_));
 sky130_fd_sc_hd__or2_1 _06914_ (.A(\_176_[5] ),
    .B(_01531_),
    .X(_01537_));
 sky130_fd_sc_hd__o211a_1 _06915_ (.A1(\_240_[5] ),
    .A2(_01526_),
    .B1(_01510_),
    .C1(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__a211o_1 _06916_ (.A1(\_243_[5] ),
    .A2(_01536_),
    .B1(_01509_),
    .C1(_01538_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _06917_ (.A0(\_176_[6] ),
    .A1(\_240_[6] ),
    .S(_01449_),
    .X(_01539_));
 sky130_fd_sc_hd__or2_1 _06918_ (.A(_01448_),
    .B(_01539_),
    .X(_01540_));
 sky130_fd_sc_hd__o211a_1 _06919_ (.A1(\_243_[6] ),
    .A2(_01485_),
    .B1(_01481_),
    .C1(_01540_),
    .X(_00185_));
 sky130_fd_sc_hd__or2_1 _06920_ (.A(\_176_[7] ),
    .B(_01531_),
    .X(_01541_));
 sky130_fd_sc_hd__o211a_1 _06921_ (.A1(\_240_[7] ),
    .A2(_01526_),
    .B1(_01510_),
    .C1(_01541_),
    .X(_01542_));
 sky130_fd_sc_hd__a211o_1 _06922_ (.A1(\_243_[7] ),
    .A2(_01536_),
    .B1(_01509_),
    .C1(_01542_),
    .X(_00186_));
 sky130_fd_sc_hd__or2_1 _06923_ (.A(\_176_[8] ),
    .B(_01531_),
    .X(_01543_));
 sky130_fd_sc_hd__o211a_1 _06924_ (.A1(\_240_[8] ),
    .A2(_01526_),
    .B1(_01510_),
    .C1(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__a211o_1 _06925_ (.A1(\_243_[8] ),
    .A2(_01536_),
    .B1(_01509_),
    .C1(_01544_),
    .X(_00187_));
 sky130_fd_sc_hd__buf_2 _06926_ (.A(_01480_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _06927_ (.A0(\_176_[9] ),
    .A1(\_240_[9] ),
    .S(_01449_),
    .X(_01546_));
 sky130_fd_sc_hd__or2_1 _06928_ (.A(_01448_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__o211a_1 _06929_ (.A1(\_243_[9] ),
    .A2(_01485_),
    .B1(_01545_),
    .C1(_01547_),
    .X(_00188_));
 sky130_fd_sc_hd__buf_2 _06930_ (.A(_01421_),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _06931_ (.A0(\_176_[10] ),
    .A1(\_240_[10] ),
    .S(_01449_),
    .X(_01549_));
 sky130_fd_sc_hd__or2_1 _06932_ (.A(_01448_),
    .B(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__o211a_1 _06933_ (.A1(\_243_[10] ),
    .A2(_01548_),
    .B1(_01545_),
    .C1(_01550_),
    .X(_00189_));
 sky130_fd_sc_hd__or2_1 _06934_ (.A(\_176_[11] ),
    .B(_01531_),
    .X(_01551_));
 sky130_fd_sc_hd__o211a_1 _06935_ (.A1(\_240_[11] ),
    .A2(_01526_),
    .B1(_01510_),
    .C1(_01551_),
    .X(_01552_));
 sky130_fd_sc_hd__a211o_1 _06936_ (.A1(\_243_[11] ),
    .A2(_01536_),
    .B1(_01509_),
    .C1(_01552_),
    .X(_00190_));
 sky130_fd_sc_hd__or2_1 _06937_ (.A(\_176_[12] ),
    .B(_01531_),
    .X(_01553_));
 sky130_fd_sc_hd__o211a_1 _06938_ (.A1(\_240_[12] ),
    .A2(_01526_),
    .B1(_01510_),
    .C1(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__a211o_1 _06939_ (.A1(\_243_[12] ),
    .A2(_01536_),
    .B1(_01509_),
    .C1(_01554_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _06940_ (.A0(\_176_[13] ),
    .A1(\_240_[13] ),
    .S(_01449_),
    .X(_01555_));
 sky130_fd_sc_hd__or2_1 _06941_ (.A(_01448_),
    .B(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__o211a_1 _06942_ (.A1(\_243_[13] ),
    .A2(_01548_),
    .B1(_01545_),
    .C1(_01556_),
    .X(_00192_));
 sky130_fd_sc_hd__clkbuf_4 _06943_ (.A(_01435_),
    .X(_01557_));
 sky130_fd_sc_hd__clkbuf_4 _06944_ (.A(_01420_),
    .X(_01558_));
 sky130_fd_sc_hd__or2_1 _06945_ (.A(\_176_[14] ),
    .B(_01531_),
    .X(_01559_));
 sky130_fd_sc_hd__o211a_1 _06946_ (.A1(\_240_[14] ),
    .A2(_01526_),
    .B1(_01558_),
    .C1(_01559_),
    .X(_01560_));
 sky130_fd_sc_hd__a211o_1 _06947_ (.A1(\_243_[14] ),
    .A2(_01536_),
    .B1(_01557_),
    .C1(_01560_),
    .X(_00193_));
 sky130_fd_sc_hd__or2_1 _06948_ (.A(\_176_[15] ),
    .B(_01531_),
    .X(_01561_));
 sky130_fd_sc_hd__o211a_1 _06949_ (.A1(\_240_[15] ),
    .A2(_01526_),
    .B1(_01558_),
    .C1(_01561_),
    .X(_01562_));
 sky130_fd_sc_hd__a211o_1 _06950_ (.A1(\_243_[15] ),
    .A2(_01536_),
    .B1(_01557_),
    .C1(_01562_),
    .X(_00194_));
 sky130_fd_sc_hd__or2_1 _06951_ (.A(\_176_[16] ),
    .B(_01531_),
    .X(_01563_));
 sky130_fd_sc_hd__o211a_1 _06952_ (.A1(\_240_[16] ),
    .A2(_01526_),
    .B1(_01558_),
    .C1(_01563_),
    .X(_01564_));
 sky130_fd_sc_hd__a211o_1 _06953_ (.A1(\_243_[16] ),
    .A2(_01536_),
    .B1(_01557_),
    .C1(_01564_),
    .X(_00195_));
 sky130_fd_sc_hd__buf_2 _06954_ (.A(_01427_),
    .X(_01565_));
 sky130_fd_sc_hd__or2_1 _06955_ (.A(\_176_[17] ),
    .B(_01531_),
    .X(_01566_));
 sky130_fd_sc_hd__o211a_1 _06956_ (.A1(\_240_[17] ),
    .A2(_01565_),
    .B1(_01558_),
    .C1(_01566_),
    .X(_01567_));
 sky130_fd_sc_hd__a211o_1 _06957_ (.A1(\_243_[17] ),
    .A2(_01536_),
    .B1(_01557_),
    .C1(_01567_),
    .X(_00196_));
 sky130_fd_sc_hd__clkbuf_2 _06958_ (.A(_01405_),
    .X(_01568_));
 sky130_fd_sc_hd__buf_4 _06959_ (.A(_01518_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _06960_ (.A0(\_176_[18] ),
    .A1(\_240_[18] ),
    .S(_01569_),
    .X(_01570_));
 sky130_fd_sc_hd__or2_1 _06961_ (.A(_01568_),
    .B(_01570_),
    .X(_01571_));
 sky130_fd_sc_hd__o211a_1 _06962_ (.A1(\_243_[18] ),
    .A2(_01548_),
    .B1(_01545_),
    .C1(_01571_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _06963_ (.A0(\_176_[19] ),
    .A1(\_240_[19] ),
    .S(_01569_),
    .X(_01572_));
 sky130_fd_sc_hd__or2_1 _06964_ (.A(_01568_),
    .B(_01572_),
    .X(_01573_));
 sky130_fd_sc_hd__o211a_1 _06965_ (.A1(\_243_[19] ),
    .A2(_01548_),
    .B1(_01545_),
    .C1(_01573_),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _06966_ (.A0(\_176_[20] ),
    .A1(\_240_[20] ),
    .S(_01569_),
    .X(_01574_));
 sky130_fd_sc_hd__or2_1 _06967_ (.A(_01568_),
    .B(_01574_),
    .X(_01575_));
 sky130_fd_sc_hd__o211a_1 _06968_ (.A1(\_243_[20] ),
    .A2(_01548_),
    .B1(_01545_),
    .C1(_01575_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _06969_ (.A0(\_176_[21] ),
    .A1(\_240_[21] ),
    .S(_01569_),
    .X(_01576_));
 sky130_fd_sc_hd__or2_1 _06970_ (.A(_01568_),
    .B(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__o211a_1 _06971_ (.A1(\_243_[21] ),
    .A2(_01548_),
    .B1(_01545_),
    .C1(_01577_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _06972_ (.A0(\_176_[22] ),
    .A1(\_240_[22] ),
    .S(_01569_),
    .X(_01578_));
 sky130_fd_sc_hd__or2_1 _06973_ (.A(_01568_),
    .B(_01578_),
    .X(_01579_));
 sky130_fd_sc_hd__o211a_1 _06974_ (.A1(\_243_[22] ),
    .A2(_01548_),
    .B1(_01545_),
    .C1(_01579_),
    .X(_00201_));
 sky130_fd_sc_hd__clkbuf_2 _06975_ (.A(_01339_),
    .X(_01580_));
 sky130_fd_sc_hd__or2_1 _06976_ (.A(\_176_[23] ),
    .B(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__o211a_1 _06977_ (.A1(\_240_[23] ),
    .A2(_01565_),
    .B1(_01558_),
    .C1(_01581_),
    .X(_01582_));
 sky130_fd_sc_hd__a211o_1 _06978_ (.A1(\_243_[23] ),
    .A2(_01536_),
    .B1(_01557_),
    .C1(_01582_),
    .X(_00202_));
 sky130_fd_sc_hd__buf_2 _06979_ (.A(_01495_),
    .X(_01583_));
 sky130_fd_sc_hd__or2_1 _06980_ (.A(\_176_[24] ),
    .B(_01580_),
    .X(_01584_));
 sky130_fd_sc_hd__o211a_1 _06981_ (.A1(\_240_[24] ),
    .A2(_01565_),
    .B1(_01558_),
    .C1(_01584_),
    .X(_01585_));
 sky130_fd_sc_hd__a211o_1 _06982_ (.A1(\_243_[24] ),
    .A2(_01583_),
    .B1(_01557_),
    .C1(_01585_),
    .X(_00203_));
 sky130_fd_sc_hd__or2_1 _06983_ (.A(\_176_[25] ),
    .B(_01580_),
    .X(_01586_));
 sky130_fd_sc_hd__o211a_1 _06984_ (.A1(\_240_[25] ),
    .A2(_01565_),
    .B1(_01558_),
    .C1(_01586_),
    .X(_01587_));
 sky130_fd_sc_hd__a211o_1 _06985_ (.A1(\_243_[25] ),
    .A2(_01583_),
    .B1(_01557_),
    .C1(_01587_),
    .X(_00204_));
 sky130_fd_sc_hd__or2_1 _06986_ (.A(\_176_[26] ),
    .B(_01580_),
    .X(_01588_));
 sky130_fd_sc_hd__o211a_1 _06987_ (.A1(\_240_[26] ),
    .A2(_01565_),
    .B1(_01558_),
    .C1(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__a211o_1 _06988_ (.A1(\_243_[26] ),
    .A2(_01583_),
    .B1(_01557_),
    .C1(_01589_),
    .X(_00205_));
 sky130_fd_sc_hd__or2_1 _06989_ (.A(\_176_[27] ),
    .B(_01580_),
    .X(_01590_));
 sky130_fd_sc_hd__o211a_1 _06990_ (.A1(\_240_[27] ),
    .A2(_01565_),
    .B1(_01558_),
    .C1(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__a211o_1 _06991_ (.A1(\_243_[27] ),
    .A2(_01583_),
    .B1(_01557_),
    .C1(_01591_),
    .X(_00206_));
 sky130_fd_sc_hd__or2_1 _06992_ (.A(\_176_[28] ),
    .B(_01580_),
    .X(_01592_));
 sky130_fd_sc_hd__o211a_1 _06993_ (.A1(\_240_[28] ),
    .A2(_01565_),
    .B1(_01558_),
    .C1(_01592_),
    .X(_01593_));
 sky130_fd_sc_hd__a211o_1 _06994_ (.A1(\_243_[28] ),
    .A2(_01583_),
    .B1(_01557_),
    .C1(_01593_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _06995_ (.A0(\_176_[29] ),
    .A1(\_240_[29] ),
    .S(_01569_),
    .X(_01594_));
 sky130_fd_sc_hd__or2_1 _06996_ (.A(_01568_),
    .B(_01594_),
    .X(_01595_));
 sky130_fd_sc_hd__o211a_1 _06997_ (.A1(\_243_[29] ),
    .A2(_01548_),
    .B1(_01545_),
    .C1(_01595_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _06998_ (.A0(\_176_[30] ),
    .A1(\_240_[30] ),
    .S(_01569_),
    .X(_01596_));
 sky130_fd_sc_hd__or2_1 _06999_ (.A(_01568_),
    .B(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__o211a_1 _07000_ (.A1(\_243_[30] ),
    .A2(_01548_),
    .B1(_01545_),
    .C1(_01597_),
    .X(_00209_));
 sky130_fd_sc_hd__buf_2 _07001_ (.A(_01480_),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _07002_ (.A0(\_176_[31] ),
    .A1(\_240_[31] ),
    .S(_01569_),
    .X(_01599_));
 sky130_fd_sc_hd__or2_1 _07003_ (.A(_01568_),
    .B(_01599_),
    .X(_01600_));
 sky130_fd_sc_hd__o211a_1 _07004_ (.A1(\_243_[31] ),
    .A2(_01548_),
    .B1(_01598_),
    .C1(_01600_),
    .X(_00210_));
 sky130_fd_sc_hd__clkbuf_4 _07005_ (.A(_01421_),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _07006_ (.A0(\_173_[0] ),
    .A1(\_237_[0] ),
    .S(_01569_),
    .X(_01602_));
 sky130_fd_sc_hd__or2_1 _07007_ (.A(_01568_),
    .B(_01602_),
    .X(_01603_));
 sky130_fd_sc_hd__o211a_1 _07008_ (.A1(\_240_[0] ),
    .A2(_01601_),
    .B1(_01598_),
    .C1(_01603_),
    .X(_00211_));
 sky130_fd_sc_hd__clkbuf_4 _07009_ (.A(\_237_[1] ),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_1 _07010_ (.A0(\_173_[1] ),
    .A1(_01604_),
    .S(_01569_),
    .X(_01605_));
 sky130_fd_sc_hd__or2_1 _07011_ (.A(_01568_),
    .B(_01605_),
    .X(_01606_));
 sky130_fd_sc_hd__o211a_1 _07012_ (.A1(\_240_[1] ),
    .A2(_01601_),
    .B1(_01598_),
    .C1(_01606_),
    .X(_00212_));
 sky130_fd_sc_hd__buf_2 _07013_ (.A(_01435_),
    .X(_01607_));
 sky130_fd_sc_hd__buf_4 _07014_ (.A(\_237_[2] ),
    .X(_01608_));
 sky130_fd_sc_hd__buf_2 _07015_ (.A(_01420_),
    .X(_01609_));
 sky130_fd_sc_hd__or2_1 _07016_ (.A(\_173_[2] ),
    .B(_01580_),
    .X(_01610_));
 sky130_fd_sc_hd__o211a_1 _07017_ (.A1(_01608_),
    .A2(_01565_),
    .B1(_01609_),
    .C1(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__a211o_1 _07018_ (.A1(\_240_[2] ),
    .A2(_01583_),
    .B1(_01607_),
    .C1(_01611_),
    .X(_00213_));
 sky130_fd_sc_hd__buf_4 _07019_ (.A(\_237_[3] ),
    .X(_01612_));
 sky130_fd_sc_hd__or2_1 _07020_ (.A(\_173_[3] ),
    .B(_01580_),
    .X(_01613_));
 sky130_fd_sc_hd__o211a_1 _07021_ (.A1(_01612_),
    .A2(_01565_),
    .B1(_01609_),
    .C1(_01613_),
    .X(_01614_));
 sky130_fd_sc_hd__a211o_1 _07022_ (.A1(\_240_[3] ),
    .A2(_01583_),
    .B1(_01607_),
    .C1(_01614_),
    .X(_00214_));
 sky130_fd_sc_hd__clkbuf_2 _07023_ (.A(_01405_),
    .X(_01615_));
 sky130_fd_sc_hd__buf_4 _07024_ (.A(\_237_[4] ),
    .X(_01616_));
 sky130_fd_sc_hd__clkbuf_4 _07025_ (.A(_01518_),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _07026_ (.A0(\_173_[4] ),
    .A1(_01616_),
    .S(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__or2_1 _07027_ (.A(_01615_),
    .B(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__o211a_1 _07028_ (.A1(\_240_[4] ),
    .A2(_01601_),
    .B1(_01598_),
    .C1(_01619_),
    .X(_00215_));
 sky130_fd_sc_hd__buf_4 _07029_ (.A(\_237_[5] ),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _07030_ (.A0(\_173_[5] ),
    .A1(_01620_),
    .S(_01617_),
    .X(_01621_));
 sky130_fd_sc_hd__or2_1 _07031_ (.A(_01615_),
    .B(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__o211a_1 _07032_ (.A1(\_240_[5] ),
    .A2(_01601_),
    .B1(_01598_),
    .C1(_01622_),
    .X(_00216_));
 sky130_fd_sc_hd__clkbuf_8 _07033_ (.A(\_237_[6] ),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _07034_ (.A0(\_173_[6] ),
    .A1(_01623_),
    .S(_01617_),
    .X(_01624_));
 sky130_fd_sc_hd__or2_1 _07035_ (.A(_01615_),
    .B(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__o211a_1 _07036_ (.A1(\_240_[6] ),
    .A2(_01601_),
    .B1(_01598_),
    .C1(_01625_),
    .X(_00217_));
 sky130_fd_sc_hd__buf_6 _07037_ (.A(\_237_[7] ),
    .X(_01626_));
 sky130_fd_sc_hd__or2_1 _07038_ (.A(\_173_[7] ),
    .B(_01580_),
    .X(_01627_));
 sky130_fd_sc_hd__o211a_1 _07039_ (.A1(_01626_),
    .A2(_01565_),
    .B1(_01609_),
    .C1(_01627_),
    .X(_01628_));
 sky130_fd_sc_hd__a211o_1 _07040_ (.A1(\_240_[7] ),
    .A2(_01583_),
    .B1(_01607_),
    .C1(_01628_),
    .X(_00218_));
 sky130_fd_sc_hd__buf_6 _07041_ (.A(\_237_[8] ),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _07042_ (.A0(\_173_[8] ),
    .A1(_01629_),
    .S(_01617_),
    .X(_01630_));
 sky130_fd_sc_hd__or2_1 _07043_ (.A(_01615_),
    .B(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__o211a_1 _07044_ (.A1(\_240_[8] ),
    .A2(_01601_),
    .B1(_01598_),
    .C1(_01631_),
    .X(_00219_));
 sky130_fd_sc_hd__buf_6 _07045_ (.A(\_237_[9] ),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _07046_ (.A0(\_173_[9] ),
    .A1(_01632_),
    .S(_01617_),
    .X(_01633_));
 sky130_fd_sc_hd__or2_1 _07047_ (.A(_01615_),
    .B(_01633_),
    .X(_01634_));
 sky130_fd_sc_hd__o211a_1 _07048_ (.A1(\_240_[9] ),
    .A2(_01601_),
    .B1(_01598_),
    .C1(_01634_),
    .X(_00220_));
 sky130_fd_sc_hd__buf_4 _07049_ (.A(\_237_[10] ),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _07050_ (.A0(\_173_[10] ),
    .A1(_01635_),
    .S(_01617_),
    .X(_01636_));
 sky130_fd_sc_hd__or2_1 _07051_ (.A(_01615_),
    .B(_01636_),
    .X(_01637_));
 sky130_fd_sc_hd__o211a_1 _07052_ (.A1(\_240_[10] ),
    .A2(_01601_),
    .B1(_01598_),
    .C1(_01637_),
    .X(_00221_));
 sky130_fd_sc_hd__buf_4 _07053_ (.A(\_237_[11] ),
    .X(_01638_));
 sky130_fd_sc_hd__buf_2 _07054_ (.A(_01427_),
    .X(_01639_));
 sky130_fd_sc_hd__or2_1 _07055_ (.A(\_173_[11] ),
    .B(_01580_),
    .X(_01640_));
 sky130_fd_sc_hd__o211a_1 _07056_ (.A1(_01638_),
    .A2(_01639_),
    .B1(_01609_),
    .C1(_01640_),
    .X(_01641_));
 sky130_fd_sc_hd__a211o_1 _07057_ (.A1(\_240_[11] ),
    .A2(_01583_),
    .B1(_01607_),
    .C1(_01641_),
    .X(_00222_));
 sky130_fd_sc_hd__buf_4 _07058_ (.A(\_237_[12] ),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _07059_ (.A0(\_173_[12] ),
    .A1(_01642_),
    .S(_01617_),
    .X(_01643_));
 sky130_fd_sc_hd__or2_1 _07060_ (.A(_01615_),
    .B(_01643_),
    .X(_01644_));
 sky130_fd_sc_hd__o211a_1 _07061_ (.A1(\_240_[12] ),
    .A2(_01601_),
    .B1(_01598_),
    .C1(_01644_),
    .X(_00223_));
 sky130_fd_sc_hd__buf_6 _07062_ (.A(\_237_[13] ),
    .X(_01645_));
 sky130_fd_sc_hd__clkbuf_2 _07063_ (.A(_01339_),
    .X(_01646_));
 sky130_fd_sc_hd__or2_1 _07064_ (.A(\_173_[13] ),
    .B(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__o211a_1 _07065_ (.A1(_01645_),
    .A2(_01639_),
    .B1(_01609_),
    .C1(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__a211o_1 _07066_ (.A1(\_240_[13] ),
    .A2(_01583_),
    .B1(_01607_),
    .C1(_01648_),
    .X(_00224_));
 sky130_fd_sc_hd__clkbuf_4 _07067_ (.A(_01495_),
    .X(_01649_));
 sky130_fd_sc_hd__buf_4 _07068_ (.A(\_237_[14] ),
    .X(_01650_));
 sky130_fd_sc_hd__or2_1 _07069_ (.A(\_173_[14] ),
    .B(_01646_),
    .X(_01651_));
 sky130_fd_sc_hd__o211a_1 _07070_ (.A1(_01650_),
    .A2(_01639_),
    .B1(_01609_),
    .C1(_01651_),
    .X(_01652_));
 sky130_fd_sc_hd__a211o_1 _07071_ (.A1(\_240_[14] ),
    .A2(_01649_),
    .B1(_01607_),
    .C1(_01652_),
    .X(_00225_));
 sky130_fd_sc_hd__clkbuf_4 _07072_ (.A(_01480_),
    .X(_01653_));
 sky130_fd_sc_hd__clkbuf_4 _07073_ (.A(\_237_[15] ),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _07074_ (.A0(\_173_[15] ),
    .A1(_01654_),
    .S(_01617_),
    .X(_01655_));
 sky130_fd_sc_hd__or2_1 _07075_ (.A(_01615_),
    .B(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__o211a_1 _07076_ (.A1(\_240_[15] ),
    .A2(_01601_),
    .B1(_01653_),
    .C1(_01656_),
    .X(_00226_));
 sky130_fd_sc_hd__buf_4 _07077_ (.A(\_237_[16] ),
    .X(_01657_));
 sky130_fd_sc_hd__or2_1 _07078_ (.A(\_173_[16] ),
    .B(_01646_),
    .X(_01658_));
 sky130_fd_sc_hd__o211a_1 _07079_ (.A1(_01657_),
    .A2(_01639_),
    .B1(_01609_),
    .C1(_01658_),
    .X(_01659_));
 sky130_fd_sc_hd__a211o_1 _07080_ (.A1(\_240_[16] ),
    .A2(_01649_),
    .B1(_01607_),
    .C1(_01659_),
    .X(_00227_));
 sky130_fd_sc_hd__buf_4 _07081_ (.A(_01421_),
    .X(_01660_));
 sky130_fd_sc_hd__clkbuf_8 _07082_ (.A(\_237_[17] ),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _07083_ (.A0(\_173_[17] ),
    .A1(_01661_),
    .S(_01617_),
    .X(_01662_));
 sky130_fd_sc_hd__or2_1 _07084_ (.A(_01615_),
    .B(_01662_),
    .X(_01663_));
 sky130_fd_sc_hd__o211a_1 _07085_ (.A1(\_240_[17] ),
    .A2(_01660_),
    .B1(_01653_),
    .C1(_01663_),
    .X(_00228_));
 sky130_fd_sc_hd__clkbuf_8 _07086_ (.A(\_237_[18] ),
    .X(_01664_));
 sky130_fd_sc_hd__or2_1 _07087_ (.A(\_173_[18] ),
    .B(_01646_),
    .X(_01665_));
 sky130_fd_sc_hd__o211a_1 _07088_ (.A1(_01664_),
    .A2(_01639_),
    .B1(_01609_),
    .C1(_01665_),
    .X(_01666_));
 sky130_fd_sc_hd__a211o_1 _07089_ (.A1(\_240_[18] ),
    .A2(_01649_),
    .B1(_01607_),
    .C1(_01666_),
    .X(_00229_));
 sky130_fd_sc_hd__buf_6 _07090_ (.A(\_237_[19] ),
    .X(_01667_));
 sky130_fd_sc_hd__mux2_1 _07091_ (.A0(\_173_[19] ),
    .A1(_01667_),
    .S(_01617_),
    .X(_01668_));
 sky130_fd_sc_hd__or2_1 _07092_ (.A(_01615_),
    .B(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__o211a_1 _07093_ (.A1(\_240_[19] ),
    .A2(_01660_),
    .B1(_01653_),
    .C1(_01669_),
    .X(_00230_));
 sky130_fd_sc_hd__buf_2 _07094_ (.A(_01405_),
    .X(_01670_));
 sky130_fd_sc_hd__buf_6 _07095_ (.A(\_237_[20] ),
    .X(_01671_));
 sky130_fd_sc_hd__buf_4 _07096_ (.A(_01518_),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _07097_ (.A0(\_173_[20] ),
    .A1(_01671_),
    .S(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__or2_1 _07098_ (.A(_01670_),
    .B(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__o211a_1 _07099_ (.A1(\_240_[20] ),
    .A2(_01660_),
    .B1(_01653_),
    .C1(_01674_),
    .X(_00231_));
 sky130_fd_sc_hd__buf_6 _07100_ (.A(\_237_[21] ),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _07101_ (.A0(\_173_[21] ),
    .A1(_01675_),
    .S(_01672_),
    .X(_01676_));
 sky130_fd_sc_hd__or2_1 _07102_ (.A(_01670_),
    .B(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__o211a_1 _07103_ (.A1(\_240_[21] ),
    .A2(_01660_),
    .B1(_01653_),
    .C1(_01677_),
    .X(_00232_));
 sky130_fd_sc_hd__buf_6 _07104_ (.A(\_237_[22] ),
    .X(_01678_));
 sky130_fd_sc_hd__mux2_1 _07105_ (.A0(\_173_[22] ),
    .A1(_01678_),
    .S(_01672_),
    .X(_01679_));
 sky130_fd_sc_hd__or2_1 _07106_ (.A(_01670_),
    .B(_01679_),
    .X(_01680_));
 sky130_fd_sc_hd__o211a_1 _07107_ (.A1(\_240_[22] ),
    .A2(_01660_),
    .B1(_01653_),
    .C1(_01680_),
    .X(_00233_));
 sky130_fd_sc_hd__buf_6 _07108_ (.A(\_237_[23] ),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _07109_ (.A0(\_173_[23] ),
    .A1(_01681_),
    .S(_01672_),
    .X(_01682_));
 sky130_fd_sc_hd__or2_1 _07110_ (.A(_01670_),
    .B(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__o211a_1 _07111_ (.A1(\_240_[23] ),
    .A2(_01660_),
    .B1(_01653_),
    .C1(_01683_),
    .X(_00234_));
 sky130_fd_sc_hd__buf_4 _07112_ (.A(\_237_[24] ),
    .X(_01684_));
 sky130_fd_sc_hd__or2_1 _07113_ (.A(\_173_[24] ),
    .B(_01646_),
    .X(_01685_));
 sky130_fd_sc_hd__o211a_1 _07114_ (.A1(_01684_),
    .A2(_01639_),
    .B1(_01609_),
    .C1(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__a211o_1 _07115_ (.A1(\_240_[24] ),
    .A2(_01649_),
    .B1(_01607_),
    .C1(_01686_),
    .X(_00235_));
 sky130_fd_sc_hd__buf_4 _07116_ (.A(\_237_[25] ),
    .X(_01687_));
 sky130_fd_sc_hd__or2_1 _07117_ (.A(\_173_[25] ),
    .B(_01646_),
    .X(_01688_));
 sky130_fd_sc_hd__o211a_1 _07118_ (.A1(_01687_),
    .A2(_01639_),
    .B1(_01609_),
    .C1(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__a211o_1 _07119_ (.A1(\_240_[25] ),
    .A2(_01649_),
    .B1(_01607_),
    .C1(_01689_),
    .X(_00236_));
 sky130_fd_sc_hd__buf_4 _07120_ (.A(\_237_[26] ),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_1 _07121_ (.A0(\_173_[26] ),
    .A1(_01690_),
    .S(_01672_),
    .X(_01691_));
 sky130_fd_sc_hd__or2_1 _07122_ (.A(_01670_),
    .B(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__o211a_1 _07123_ (.A1(\_240_[26] ),
    .A2(_01660_),
    .B1(_01653_),
    .C1(_01692_),
    .X(_00237_));
 sky130_fd_sc_hd__clkbuf_4 _07124_ (.A(_01435_),
    .X(_01693_));
 sky130_fd_sc_hd__buf_4 _07125_ (.A(\_237_[27] ),
    .X(_01694_));
 sky130_fd_sc_hd__clkbuf_4 _07126_ (.A(_01420_),
    .X(_01695_));
 sky130_fd_sc_hd__or2_1 _07127_ (.A(\_173_[27] ),
    .B(_01646_),
    .X(_01696_));
 sky130_fd_sc_hd__o211a_1 _07128_ (.A1(_01694_),
    .A2(_01639_),
    .B1(_01695_),
    .C1(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__a211o_1 _07129_ (.A1(\_240_[27] ),
    .A2(_01649_),
    .B1(_01693_),
    .C1(_01697_),
    .X(_00238_));
 sky130_fd_sc_hd__clkbuf_8 _07130_ (.A(\_237_[28] ),
    .X(_01698_));
 sky130_fd_sc_hd__or2_1 _07131_ (.A(\_173_[28] ),
    .B(_01646_),
    .X(_01699_));
 sky130_fd_sc_hd__o211a_1 _07132_ (.A1(_01698_),
    .A2(_01639_),
    .B1(_01695_),
    .C1(_01699_),
    .X(_01700_));
 sky130_fd_sc_hd__a211o_1 _07133_ (.A1(\_240_[28] ),
    .A2(_01649_),
    .B1(_01693_),
    .C1(_01700_),
    .X(_00239_));
 sky130_fd_sc_hd__buf_6 _07134_ (.A(\_237_[29] ),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _07135_ (.A0(\_173_[29] ),
    .A1(_01701_),
    .S(_01672_),
    .X(_01702_));
 sky130_fd_sc_hd__or2_1 _07136_ (.A(_01670_),
    .B(_01702_),
    .X(_01703_));
 sky130_fd_sc_hd__o211a_1 _07137_ (.A1(\_240_[29] ),
    .A2(_01660_),
    .B1(_01653_),
    .C1(_01703_),
    .X(_00240_));
 sky130_fd_sc_hd__buf_6 _07138_ (.A(\_237_[30] ),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _07139_ (.A0(\_173_[30] ),
    .A1(_01704_),
    .S(_01672_),
    .X(_01705_));
 sky130_fd_sc_hd__or2_1 _07140_ (.A(_01670_),
    .B(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__o211a_1 _07141_ (.A1(\_240_[30] ),
    .A2(_01660_),
    .B1(_01653_),
    .C1(_01706_),
    .X(_00241_));
 sky130_fd_sc_hd__buf_6 _07142_ (.A(\_237_[31] ),
    .X(_01707_));
 sky130_fd_sc_hd__or2_1 _07143_ (.A(\_173_[31] ),
    .B(_01646_),
    .X(_01708_));
 sky130_fd_sc_hd__o211a_1 _07144_ (.A1(_01707_),
    .A2(_01639_),
    .B1(_01695_),
    .C1(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__a211o_1 _07145_ (.A1(\_240_[31] ),
    .A2(_01649_),
    .B1(_01693_),
    .C1(_01709_),
    .X(_00242_));
 sky130_fd_sc_hd__buf_4 _07146_ (.A(_01417_),
    .X(_01710_));
 sky130_fd_sc_hd__nand2_2 _07147_ (.A(\_182_[0] ),
    .B(\_237_[0] ),
    .Y(_01711_));
 sky130_fd_sc_hd__or2_1 _07148_ (.A(\_182_[0] ),
    .B(\_237_[0] ),
    .X(_01712_));
 sky130_fd_sc_hd__xnor2_1 _07149_ (.A(_01638_),
    .B(_01623_),
    .Y(_01713_));
 sky130_fd_sc_hd__xnor2_2 _07150_ (.A(_01687_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__nand2_1 _07151_ (.A(\_185_[0] ),
    .B(\_234_[0] ),
    .Y(_01715_));
 sky130_fd_sc_hd__or2_1 _07152_ (.A(\_185_[0] ),
    .B(\_234_[0] ),
    .X(_01716_));
 sky130_fd_sc_hd__nand2_1 _07153_ (.A(_01715_),
    .B(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__xnor2_1 _07154_ (.A(_01714_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__mux2_1 _07155_ (.A0(\_243_[0] ),
    .A1(\_240_[0] ),
    .S(\_237_[0] ),
    .X(_01719_));
 sky130_fd_sc_hd__and2_1 _07156_ (.A(_01718_),
    .B(_01719_),
    .X(_01720_));
 sky130_fd_sc_hd__o21ai_1 _07157_ (.A1(_01718_),
    .A2(_01719_),
    .B1(_01302_),
    .Y(_01721_));
 sky130_fd_sc_hd__nor2_1 _07158_ (.A(_01720_),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__a31o_1 _07159_ (.A1(_01269_),
    .A2(_01711_),
    .A3(_01712_),
    .B1(_01722_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _07160_ (.A0(\_237_[0] ),
    .A1(_01723_),
    .S(_01411_),
    .X(_01724_));
 sky130_fd_sc_hd__or2_1 _07161_ (.A(_01710_),
    .B(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__clkbuf_1 _07162_ (.A(_01725_),
    .X(_00243_));
 sky130_fd_sc_hd__xnor2_1 _07163_ (.A(_01642_),
    .B(_01626_),
    .Y(_01726_));
 sky130_fd_sc_hd__xnor2_2 _07164_ (.A(_01690_),
    .B(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__and2_1 _07165_ (.A(\_185_[1] ),
    .B(\_234_[1] ),
    .X(_01728_));
 sky130_fd_sc_hd__nor2_1 _07166_ (.A(\_185_[1] ),
    .B(\_234_[1] ),
    .Y(_01729_));
 sky130_fd_sc_hd__nor2_1 _07167_ (.A(_01728_),
    .B(_01729_),
    .Y(_01730_));
 sky130_fd_sc_hd__xnor2_1 _07168_ (.A(_01727_),
    .B(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__a21boi_1 _07169_ (.A1(_01714_),
    .A2(_01716_),
    .B1_N(_01715_),
    .Y(_01732_));
 sky130_fd_sc_hd__xnor2_1 _07170_ (.A(_01731_),
    .B(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__mux2_2 _07171_ (.A0(\_243_[1] ),
    .A1(\_240_[1] ),
    .S(_01604_),
    .X(_01734_));
 sky130_fd_sc_hd__xnor2_1 _07172_ (.A(_01733_),
    .B(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__and2_1 _07173_ (.A(_01720_),
    .B(_01735_),
    .X(_01736_));
 sky130_fd_sc_hd__o21ai_1 _07174_ (.A1(_01720_),
    .A2(_01735_),
    .B1(_01518_),
    .Y(_01737_));
 sky130_fd_sc_hd__and2_1 _07175_ (.A(\_182_[1] ),
    .B(_01604_),
    .X(_01738_));
 sky130_fd_sc_hd__nor2_1 _07176_ (.A(\_182_[1] ),
    .B(_01604_),
    .Y(_01739_));
 sky130_fd_sc_hd__nor2_1 _07177_ (.A(_01738_),
    .B(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__xnor2_1 _07178_ (.A(_01711_),
    .B(_01740_),
    .Y(_01741_));
 sky130_fd_sc_hd__a2bb2o_1 _07179_ (.A1_N(_01736_),
    .A2_N(_01737_),
    .B1(_01269_),
    .B2(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__mux2_1 _07180_ (.A0(_01604_),
    .A1(_01742_),
    .S(_01411_),
    .X(_01743_));
 sky130_fd_sc_hd__or2_1 _07181_ (.A(_01710_),
    .B(_01743_),
    .X(_01744_));
 sky130_fd_sc_hd__clkbuf_1 _07182_ (.A(_01744_),
    .X(_00244_));
 sky130_fd_sc_hd__nand2_1 _07183_ (.A(\_182_[1] ),
    .B(_01604_),
    .Y(_01745_));
 sky130_fd_sc_hd__o21a_1 _07184_ (.A1(_01711_),
    .A2(_01739_),
    .B1(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__nand2_1 _07185_ (.A(\_182_[2] ),
    .B(_01608_),
    .Y(_01747_));
 sky130_fd_sc_hd__inv_2 _07186_ (.A(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_1 _07187_ (.A(\_182_[2] ),
    .B(_01608_),
    .Y(_01749_));
 sky130_fd_sc_hd__nor2_1 _07188_ (.A(_01748_),
    .B(_01749_),
    .Y(_01750_));
 sky130_fd_sc_hd__xnor2_1 _07189_ (.A(_01746_),
    .B(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__nor2_1 _07190_ (.A(_01731_),
    .B(_01732_),
    .Y(_01752_));
 sky130_fd_sc_hd__and2b_1 _07191_ (.A_N(_01733_),
    .B(_01734_),
    .X(_01753_));
 sky130_fd_sc_hd__xnor2_1 _07192_ (.A(_01645_),
    .B(_01629_),
    .Y(_01754_));
 sky130_fd_sc_hd__xnor2_2 _07193_ (.A(_01694_),
    .B(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__nand2_1 _07194_ (.A(\_185_[2] ),
    .B(\_234_[2] ),
    .Y(_01756_));
 sky130_fd_sc_hd__or2_1 _07195_ (.A(\_185_[2] ),
    .B(\_234_[2] ),
    .X(_01757_));
 sky130_fd_sc_hd__nand2_1 _07196_ (.A(_01756_),
    .B(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__xor2_1 _07197_ (.A(_01755_),
    .B(_01758_),
    .X(_01759_));
 sky130_fd_sc_hd__a21oi_1 _07198_ (.A1(_01727_),
    .A2(_01730_),
    .B1(_01728_),
    .Y(_01760_));
 sky130_fd_sc_hd__xnor2_1 _07199_ (.A(_01759_),
    .B(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__mux2_2 _07200_ (.A0(\_243_[2] ),
    .A1(\_240_[2] ),
    .S(_01608_),
    .X(_01762_));
 sky130_fd_sc_hd__xnor2_1 _07201_ (.A(_01761_),
    .B(_01762_),
    .Y(_01763_));
 sky130_fd_sc_hd__o21ai_1 _07202_ (.A1(_01752_),
    .A2(_01753_),
    .B1(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__or3_1 _07203_ (.A(_01752_),
    .B(_01753_),
    .C(_01763_),
    .X(_01765_));
 sky130_fd_sc_hd__and3_1 _07204_ (.A(_01736_),
    .B(_01764_),
    .C(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__a21oi_1 _07205_ (.A1(_01764_),
    .A2(_01765_),
    .B1(_01736_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_1 _07206_ (.A(_01766_),
    .B(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__mux2_1 _07207_ (.A0(_01751_),
    .A1(_01768_),
    .S(_01518_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _07208_ (.A0(_01608_),
    .A1(_01769_),
    .S(_01411_),
    .X(_01770_));
 sky130_fd_sc_hd__or2_1 _07209_ (.A(_01710_),
    .B(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__clkbuf_1 _07210_ (.A(_01771_),
    .X(_00245_));
 sky130_fd_sc_hd__nor2_1 _07211_ (.A(\_182_[3] ),
    .B(_01612_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand2_1 _07212_ (.A(\_182_[3] ),
    .B(_01612_),
    .Y(_01773_));
 sky130_fd_sc_hd__or2b_1 _07213_ (.A(_01772_),
    .B_N(_01773_),
    .X(_01774_));
 sky130_fd_sc_hd__o211a_1 _07214_ (.A1(_01711_),
    .A2(_01739_),
    .B1(_01747_),
    .C1(_01745_),
    .X(_01775_));
 sky130_fd_sc_hd__nor2_1 _07215_ (.A(_01749_),
    .B(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__xnor2_1 _07216_ (.A(_01774_),
    .B(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__clkbuf_4 _07217_ (.A(_01353_),
    .X(_01778_));
 sky130_fd_sc_hd__nand3_1 _07218_ (.A(_01755_),
    .B(_01756_),
    .C(_01757_),
    .Y(_01779_));
 sky130_fd_sc_hd__xnor2_1 _07219_ (.A(_01650_),
    .B(_01632_),
    .Y(_01780_));
 sky130_fd_sc_hd__xnor2_2 _07220_ (.A(_01698_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__nand2_1 _07221_ (.A(\_185_[3] ),
    .B(\_234_[3] ),
    .Y(_01782_));
 sky130_fd_sc_hd__or2_1 _07222_ (.A(\_185_[3] ),
    .B(\_234_[3] ),
    .X(_01783_));
 sky130_fd_sc_hd__nand2_1 _07223_ (.A(_01782_),
    .B(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__xor2_1 _07224_ (.A(_01781_),
    .B(_01784_),
    .X(_01785_));
 sky130_fd_sc_hd__a21oi_1 _07225_ (.A1(_01756_),
    .A2(_01779_),
    .B1(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__and3_1 _07226_ (.A(_01756_),
    .B(_01779_),
    .C(_01785_),
    .X(_01787_));
 sky130_fd_sc_hd__or2_1 _07227_ (.A(_01786_),
    .B(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_2 _07228_ (.A0(\_243_[3] ),
    .A1(\_240_[3] ),
    .S(_01612_),
    .X(_01789_));
 sky130_fd_sc_hd__xnor2_1 _07229_ (.A(_01788_),
    .B(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__and2b_1 _07230_ (.A_N(_01761_),
    .B(_01762_),
    .X(_01791_));
 sky130_fd_sc_hd__o21bai_1 _07231_ (.A1(_01759_),
    .A2(_01760_),
    .B1_N(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__nand2_1 _07232_ (.A(_01790_),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__or2_1 _07233_ (.A(_01790_),
    .B(_01792_),
    .X(_01794_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(_01793_),
    .B(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__a21bo_1 _07235_ (.A1(_01736_),
    .A2(_01765_),
    .B1_N(_01764_),
    .X(_01796_));
 sky130_fd_sc_hd__xor2_1 _07236_ (.A(_01795_),
    .B(_01796_),
    .X(_01797_));
 sky130_fd_sc_hd__nand2_1 _07237_ (.A(_01778_),
    .B(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__buf_4 _07238_ (.A(_01412_),
    .X(_01799_));
 sky130_fd_sc_hd__o211a_1 _07239_ (.A1(_01520_),
    .A2(_01777_),
    .B1(_01798_),
    .C1(_01799_),
    .X(_01800_));
 sky130_fd_sc_hd__a211o_1 _07240_ (.A1(_01612_),
    .A2(_01649_),
    .B1(_01693_),
    .C1(_01800_),
    .X(_00246_));
 sky130_fd_sc_hd__buf_4 _07241_ (.A(_01437_),
    .X(_01801_));
 sky130_fd_sc_hd__a21bo_1 _07242_ (.A1(_01794_),
    .A2(_01796_),
    .B1_N(_01793_),
    .X(_01802_));
 sky130_fd_sc_hd__and2b_1 _07243_ (.A_N(_01788_),
    .B(_01789_),
    .X(_01803_));
 sky130_fd_sc_hd__nand3_1 _07244_ (.A(_01781_),
    .B(_01782_),
    .C(_01783_),
    .Y(_01804_));
 sky130_fd_sc_hd__xnor2_1 _07245_ (.A(_01654_),
    .B(_01635_),
    .Y(_01805_));
 sky130_fd_sc_hd__xnor2_1 _07246_ (.A(_01701_),
    .B(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__nand2_1 _07247_ (.A(\_185_[4] ),
    .B(\_234_[4] ),
    .Y(_01807_));
 sky130_fd_sc_hd__or2_1 _07248_ (.A(\_185_[4] ),
    .B(\_234_[4] ),
    .X(_01808_));
 sky130_fd_sc_hd__nand2_1 _07249_ (.A(_01807_),
    .B(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__xor2_1 _07250_ (.A(_01806_),
    .B(_01809_),
    .X(_01810_));
 sky130_fd_sc_hd__a21oi_1 _07251_ (.A1(_01782_),
    .A2(_01804_),
    .B1(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__and3_1 _07252_ (.A(_01782_),
    .B(_01804_),
    .C(_01810_),
    .X(_01812_));
 sky130_fd_sc_hd__or2_1 _07253_ (.A(_01811_),
    .B(_01812_),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_2 _07254_ (.A0(\_243_[4] ),
    .A1(\_240_[4] ),
    .S(_01616_),
    .X(_01814_));
 sky130_fd_sc_hd__xnor2_1 _07255_ (.A(_01813_),
    .B(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__o21a_1 _07256_ (.A1(_01786_),
    .A2(_01803_),
    .B1(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__nor3_1 _07257_ (.A(_01786_),
    .B(_01803_),
    .C(_01815_),
    .Y(_01817_));
 sky130_fd_sc_hd__nor2_1 _07258_ (.A(_01816_),
    .B(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__xor2_1 _07259_ (.A(_01802_),
    .B(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__or2_1 _07260_ (.A(\_182_[4] ),
    .B(_01616_),
    .X(_01820_));
 sky130_fd_sc_hd__nand2_1 _07261_ (.A(\_182_[4] ),
    .B(_01616_),
    .Y(_01821_));
 sky130_fd_sc_hd__nand2_1 _07262_ (.A(_01820_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__o31a_2 _07263_ (.A1(_01749_),
    .A2(_01772_),
    .A3(_01775_),
    .B1(_01773_),
    .X(_01823_));
 sky130_fd_sc_hd__xnor2_2 _07264_ (.A(_01822_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__nand2_1 _07265_ (.A(_01409_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__o211a_1 _07266_ (.A1(_01801_),
    .A2(_01819_),
    .B1(_01825_),
    .C1(_01799_),
    .X(_01826_));
 sky130_fd_sc_hd__a211o_1 _07267_ (.A1(_01616_),
    .A2(_01649_),
    .B1(_01693_),
    .C1(_01826_),
    .X(_00247_));
 sky130_fd_sc_hd__clkbuf_4 _07268_ (.A(_01406_),
    .X(_01827_));
 sky130_fd_sc_hd__or2_1 _07269_ (.A(\_182_[5] ),
    .B(_01620_),
    .X(_01828_));
 sky130_fd_sc_hd__nand2_1 _07270_ (.A(\_182_[5] ),
    .B(_01620_),
    .Y(_01829_));
 sky130_fd_sc_hd__nand2_1 _07271_ (.A(_01828_),
    .B(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__o21a_1 _07272_ (.A1(_01822_),
    .A2(_01823_),
    .B1(_01821_),
    .X(_01831_));
 sky130_fd_sc_hd__xnor2_1 _07273_ (.A(_01830_),
    .B(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__inv_2 _07274_ (.A(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__and2b_1 _07275_ (.A_N(_01813_),
    .B(_01814_),
    .X(_01834_));
 sky130_fd_sc_hd__inv_2 _07276_ (.A(_01806_),
    .Y(_01835_));
 sky130_fd_sc_hd__or2_1 _07277_ (.A(_01835_),
    .B(_01809_),
    .X(_01836_));
 sky130_fd_sc_hd__xnor2_1 _07278_ (.A(_01657_),
    .B(_01638_),
    .Y(_01837_));
 sky130_fd_sc_hd__xnor2_2 _07279_ (.A(_01704_),
    .B(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__or2_1 _07280_ (.A(\_185_[5] ),
    .B(\_234_[5] ),
    .X(_01839_));
 sky130_fd_sc_hd__nand2_1 _07281_ (.A(\_185_[5] ),
    .B(\_234_[5] ),
    .Y(_01840_));
 sky130_fd_sc_hd__nand3_1 _07282_ (.A(_01838_),
    .B(_01839_),
    .C(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__a21o_1 _07283_ (.A1(_01839_),
    .A2(_01840_),
    .B1(_01838_),
    .X(_01842_));
 sky130_fd_sc_hd__nand2_1 _07284_ (.A(_01841_),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__a21oi_1 _07285_ (.A1(_01807_),
    .A2(_01836_),
    .B1(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__and3_1 _07286_ (.A(_01807_),
    .B(_01836_),
    .C(_01843_),
    .X(_01845_));
 sky130_fd_sc_hd__or2_1 _07287_ (.A(_01844_),
    .B(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_4 _07288_ (.A0(\_243_[5] ),
    .A1(\_240_[5] ),
    .S(_01620_),
    .X(_01847_));
 sky130_fd_sc_hd__xnor2_1 _07289_ (.A(_01846_),
    .B(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor3_1 _07290_ (.A(_01811_),
    .B(_01834_),
    .C(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__o21a_1 _07291_ (.A1(_01811_),
    .A2(_01834_),
    .B1(_01848_),
    .X(_01850_));
 sky130_fd_sc_hd__a21oi_1 _07292_ (.A1(_01802_),
    .A2(_01818_),
    .B1(_01816_),
    .Y(_01851_));
 sky130_fd_sc_hd__o21ai_1 _07293_ (.A1(_01849_),
    .A2(_01850_),
    .B1(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__or3_1 _07294_ (.A(_01849_),
    .B(_01850_),
    .C(_01851_),
    .X(_01853_));
 sky130_fd_sc_hd__a21o_1 _07295_ (.A1(_01852_),
    .A2(_01853_),
    .B1(_01427_),
    .X(_01854_));
 sky130_fd_sc_hd__o211a_1 _07296_ (.A1(_01520_),
    .A2(_01833_),
    .B1(_01854_),
    .C1(_01799_),
    .X(_01855_));
 sky130_fd_sc_hd__a211o_1 _07297_ (.A1(_01620_),
    .A2(_01827_),
    .B1(_01693_),
    .C1(_01855_),
    .X(_00248_));
 sky130_fd_sc_hd__clkbuf_8 _07298_ (.A(_01427_),
    .X(_01856_));
 sky130_fd_sc_hd__or2_1 _07299_ (.A(\_182_[6] ),
    .B(_01623_),
    .X(_01857_));
 sky130_fd_sc_hd__nand2_1 _07300_ (.A(\_182_[6] ),
    .B(_01623_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand2_1 _07301_ (.A(_01857_),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_1 _07302_ (.A(\_182_[5] ),
    .B(_01620_),
    .Y(_01860_));
 sky130_fd_sc_hd__nand3_1 _07303_ (.A(\_182_[4] ),
    .B(_01616_),
    .C(_01828_),
    .Y(_01861_));
 sky130_fd_sc_hd__o311a_1 _07304_ (.A1(_01822_),
    .A2(_01823_),
    .A3(_01860_),
    .B1(_01829_),
    .C1(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__xnor2_2 _07305_ (.A(_01859_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__or3_1 _07306_ (.A(_01811_),
    .B(_01834_),
    .C(_01848_),
    .X(_01864_));
 sky130_fd_sc_hd__and2b_1 _07307_ (.A_N(_01846_),
    .B(_01847_),
    .X(_01865_));
 sky130_fd_sc_hd__xnor2_1 _07308_ (.A(_01661_),
    .B(_01642_),
    .Y(_01866_));
 sky130_fd_sc_hd__xnor2_2 _07309_ (.A(_01707_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__nand2_1 _07310_ (.A(\_185_[6] ),
    .B(\_234_[6] ),
    .Y(_01868_));
 sky130_fd_sc_hd__or2_1 _07311_ (.A(\_185_[6] ),
    .B(\_234_[6] ),
    .X(_01869_));
 sky130_fd_sc_hd__nand2_1 _07312_ (.A(_01868_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__xor2_1 _07313_ (.A(_01867_),
    .B(_01870_),
    .X(_01871_));
 sky130_fd_sc_hd__a21o_1 _07314_ (.A1(_01840_),
    .A2(_01841_),
    .B1(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__nand3_1 _07315_ (.A(_01840_),
    .B(_01841_),
    .C(_01871_),
    .Y(_01873_));
 sky130_fd_sc_hd__nand2_1 _07316_ (.A(_01872_),
    .B(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__mux2_4 _07317_ (.A0(\_243_[6] ),
    .A1(\_240_[6] ),
    .S(_01623_),
    .X(_01875_));
 sky130_fd_sc_hd__xnor2_1 _07318_ (.A(_01874_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__o21a_1 _07319_ (.A1(_01844_),
    .A2(_01865_),
    .B1(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__nor3_1 _07320_ (.A(_01844_),
    .B(_01865_),
    .C(_01876_),
    .Y(_01878_));
 sky130_fd_sc_hd__nor2_1 _07321_ (.A(_01877_),
    .B(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__a211o_1 _07322_ (.A1(_01802_),
    .A2(_01818_),
    .B1(_01850_),
    .C1(_01816_),
    .X(_01880_));
 sky130_fd_sc_hd__and3_1 _07323_ (.A(_01864_),
    .B(_01879_),
    .C(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__a21oi_1 _07324_ (.A1(_01864_),
    .A2(_01880_),
    .B1(_01879_),
    .Y(_01882_));
 sky130_fd_sc_hd__o21a_1 _07325_ (.A1(_01881_),
    .A2(_01882_),
    .B1(_01354_),
    .X(_01883_));
 sky130_fd_sc_hd__clkbuf_8 _07326_ (.A(_01405_),
    .X(_01884_));
 sky130_fd_sc_hd__a211oi_1 _07327_ (.A1(_01856_),
    .A2(_01863_),
    .B1(_01883_),
    .C1(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__a211o_1 _07328_ (.A1(_01623_),
    .A2(_01827_),
    .B1(_01693_),
    .C1(_01885_),
    .X(_00249_));
 sky130_fd_sc_hd__buf_4 _07329_ (.A(_01480_),
    .X(_01886_));
 sky130_fd_sc_hd__or2_1 _07330_ (.A(\_182_[7] ),
    .B(_01626_),
    .X(_01887_));
 sky130_fd_sc_hd__nand2_1 _07331_ (.A(\_182_[7] ),
    .B(_01626_),
    .Y(_01888_));
 sky130_fd_sc_hd__nand2_1 _07332_ (.A(_01887_),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__o21a_1 _07333_ (.A1(_01859_),
    .A2(_01862_),
    .B1(_01858_),
    .X(_01890_));
 sky130_fd_sc_hd__xnor2_1 _07334_ (.A(_01889_),
    .B(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__inv_2 _07335_ (.A(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__or2b_1 _07336_ (.A(_01874_),
    .B_N(_01875_),
    .X(_01893_));
 sky130_fd_sc_hd__nand3_1 _07337_ (.A(_01867_),
    .B(_01868_),
    .C(_01869_),
    .Y(_01894_));
 sky130_fd_sc_hd__xnor2_1 _07338_ (.A(_01645_),
    .B(\_237_[0] ),
    .Y(_01895_));
 sky130_fd_sc_hd__xnor2_1 _07339_ (.A(_01664_),
    .B(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__nand2_1 _07340_ (.A(\_185_[7] ),
    .B(\_234_[7] ),
    .Y(_01897_));
 sky130_fd_sc_hd__or2_1 _07341_ (.A(\_185_[7] ),
    .B(\_234_[7] ),
    .X(_01898_));
 sky130_fd_sc_hd__nand2_1 _07342_ (.A(_01897_),
    .B(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__xor2_1 _07343_ (.A(_01896_),
    .B(_01899_),
    .X(_01900_));
 sky130_fd_sc_hd__a21oi_1 _07344_ (.A1(_01868_),
    .A2(_01894_),
    .B1(_01900_),
    .Y(_01901_));
 sky130_fd_sc_hd__and3_1 _07345_ (.A(_01868_),
    .B(_01894_),
    .C(_01900_),
    .X(_01902_));
 sky130_fd_sc_hd__or2_1 _07346_ (.A(_01901_),
    .B(_01902_),
    .X(_01903_));
 sky130_fd_sc_hd__nor2_1 _07347_ (.A(_01626_),
    .B(\_243_[7] ),
    .Y(_01904_));
 sky130_fd_sc_hd__and2b_1 _07348_ (.A_N(\_240_[7] ),
    .B(_01626_),
    .X(_01905_));
 sky130_fd_sc_hd__nor2_2 _07349_ (.A(_01904_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__xor2_1 _07350_ (.A(_01903_),
    .B(_01906_),
    .X(_01907_));
 sky130_fd_sc_hd__a21oi_1 _07351_ (.A1(_01872_),
    .A2(_01893_),
    .B1(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__nand3_1 _07352_ (.A(_01872_),
    .B(_01893_),
    .C(_01907_),
    .Y(_01909_));
 sky130_fd_sc_hd__or2b_1 _07353_ (.A(_01908_),
    .B_N(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__inv_2 _07354_ (.A(_01910_),
    .Y(_01911_));
 sky130_fd_sc_hd__or2_1 _07355_ (.A(_01877_),
    .B(_01881_),
    .X(_01912_));
 sky130_fd_sc_hd__o21ai_1 _07356_ (.A1(_01911_),
    .A2(_01912_),
    .B1(_01523_),
    .Y(_01913_));
 sky130_fd_sc_hd__a21oi_1 _07357_ (.A1(_01911_),
    .A2(_01912_),
    .B1(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__a211o_1 _07358_ (.A1(_01856_),
    .A2(_01892_),
    .B1(_01914_),
    .C1(_01884_),
    .X(_01915_));
 sky130_fd_sc_hd__o211a_1 _07359_ (.A1(_01626_),
    .A2(_01660_),
    .B1(_01886_),
    .C1(_01915_),
    .X(_00250_));
 sky130_fd_sc_hd__or2_1 _07360_ (.A(\_182_[8] ),
    .B(_01629_),
    .X(_01916_));
 sky130_fd_sc_hd__nand2_1 _07361_ (.A(\_182_[8] ),
    .B(_01629_),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_2 _07362_ (.A(_01916_),
    .B(_01917_),
    .Y(_01918_));
 sky130_fd_sc_hd__and3_1 _07363_ (.A(\_182_[6] ),
    .B(_01623_),
    .C(_01887_),
    .X(_01919_));
 sky130_fd_sc_hd__a21oi_1 _07364_ (.A1(\_182_[7] ),
    .A2(_01626_),
    .B1(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hd__o31a_2 _07365_ (.A1(_01859_),
    .A2(_01862_),
    .A3(_01889_),
    .B1(_01920_),
    .X(_01921_));
 sky130_fd_sc_hd__xnor2_4 _07366_ (.A(_01918_),
    .B(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__clkbuf_8 _07367_ (.A(_01408_),
    .X(_01923_));
 sky130_fd_sc_hd__o21a_1 _07368_ (.A1(_01877_),
    .A2(_01908_),
    .B1(_01909_),
    .X(_01924_));
 sky130_fd_sc_hd__and4_1 _07369_ (.A(_01864_),
    .B(_01879_),
    .C(_01880_),
    .D(_01911_),
    .X(_01925_));
 sky130_fd_sc_hd__and2b_1 _07370_ (.A_N(_01903_),
    .B(_01906_),
    .X(_01926_));
 sky130_fd_sc_hd__inv_2 _07371_ (.A(_01896_),
    .Y(_01927_));
 sky130_fd_sc_hd__or2_1 _07372_ (.A(_01927_),
    .B(_01899_),
    .X(_01928_));
 sky130_fd_sc_hd__xnor2_1 _07373_ (.A(_01650_),
    .B(_01604_),
    .Y(_01929_));
 sky130_fd_sc_hd__xnor2_2 _07374_ (.A(_01667_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__or2_1 _07375_ (.A(\_185_[8] ),
    .B(\_234_[8] ),
    .X(_01931_));
 sky130_fd_sc_hd__nand2_1 _07376_ (.A(\_185_[8] ),
    .B(\_234_[8] ),
    .Y(_01932_));
 sky130_fd_sc_hd__nand3_1 _07377_ (.A(_01930_),
    .B(_01931_),
    .C(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__a21o_1 _07378_ (.A1(_01931_),
    .A2(_01932_),
    .B1(_01930_),
    .X(_01934_));
 sky130_fd_sc_hd__nand2_1 _07379_ (.A(_01933_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__a21oi_1 _07380_ (.A1(_01897_),
    .A2(_01928_),
    .B1(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__and3_1 _07381_ (.A(_01897_),
    .B(_01928_),
    .C(_01935_),
    .X(_01937_));
 sky130_fd_sc_hd__or2_1 _07382_ (.A(_01936_),
    .B(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_4 _07383_ (.A0(\_243_[8] ),
    .A1(\_240_[8] ),
    .S(_01629_),
    .X(_01939_));
 sky130_fd_sc_hd__xnor2_1 _07384_ (.A(_01938_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__o21a_1 _07385_ (.A1(_01901_),
    .A2(_01926_),
    .B1(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__nor3_1 _07386_ (.A(_01901_),
    .B(_01926_),
    .C(_01940_),
    .Y(_01942_));
 sky130_fd_sc_hd__nor2_1 _07387_ (.A(_01941_),
    .B(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__o21a_1 _07388_ (.A1(_01924_),
    .A2(_01925_),
    .B1(_01943_),
    .X(_01944_));
 sky130_fd_sc_hd__nor2_1 _07389_ (.A(_01923_),
    .B(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__or3_1 _07390_ (.A(_01943_),
    .B(_01924_),
    .C(_01925_),
    .X(_01946_));
 sky130_fd_sc_hd__a2bb2o_1 _07391_ (.A1_N(_01520_),
    .A2_N(_01922_),
    .B1(_01945_),
    .B2(_01946_),
    .X(_01947_));
 sky130_fd_sc_hd__or2_1 _07392_ (.A(_01629_),
    .B(_01412_),
    .X(_01948_));
 sky130_fd_sc_hd__buf_4 _07393_ (.A(_01480_),
    .X(_00105_));
 sky130_fd_sc_hd__o211a_1 _07394_ (.A1(_01407_),
    .A2(_01947_),
    .B1(_01948_),
    .C1(_00105_),
    .X(_00251_));
 sky130_fd_sc_hd__nor2_1 _07395_ (.A(_01941_),
    .B(_01944_),
    .Y(_01949_));
 sky130_fd_sc_hd__and2b_1 _07396_ (.A_N(_01938_),
    .B(_01939_),
    .X(_01950_));
 sky130_fd_sc_hd__xnor2_1 _07397_ (.A(_01654_),
    .B(_01608_),
    .Y(_01951_));
 sky130_fd_sc_hd__xnor2_1 _07398_ (.A(_01671_),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__or2_1 _07399_ (.A(\_185_[9] ),
    .B(\_234_[9] ),
    .X(_01953_));
 sky130_fd_sc_hd__nand2_1 _07400_ (.A(\_185_[9] ),
    .B(\_234_[9] ),
    .Y(_01954_));
 sky130_fd_sc_hd__nand2_1 _07401_ (.A(_01953_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__xor2_1 _07402_ (.A(_01952_),
    .B(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__a21oi_1 _07403_ (.A1(_01932_),
    .A2(_01933_),
    .B1(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__and3_1 _07404_ (.A(_01932_),
    .B(_01933_),
    .C(_01956_),
    .X(_01958_));
 sky130_fd_sc_hd__or2_1 _07405_ (.A(_01957_),
    .B(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_2 _07406_ (.A0(\_243_[9] ),
    .A1(\_240_[9] ),
    .S(_01632_),
    .X(_01960_));
 sky130_fd_sc_hd__xnor2_1 _07407_ (.A(_01959_),
    .B(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__or3_1 _07408_ (.A(_01936_),
    .B(_01950_),
    .C(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__o21ai_1 _07409_ (.A1(_01936_),
    .A2(_01950_),
    .B1(_01961_),
    .Y(_01963_));
 sky130_fd_sc_hd__and2_1 _07410_ (.A(_01962_),
    .B(_01963_),
    .X(_01964_));
 sky130_fd_sc_hd__nand2_1 _07411_ (.A(_01949_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__o21a_1 _07412_ (.A1(_01949_),
    .A2(_01964_),
    .B1(_01354_),
    .X(_01966_));
 sky130_fd_sc_hd__or2_1 _07413_ (.A(\_182_[9] ),
    .B(_01632_),
    .X(_01967_));
 sky130_fd_sc_hd__nand2_1 _07414_ (.A(\_182_[9] ),
    .B(_01632_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_2 _07415_ (.A(_01967_),
    .B(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__o21ai_2 _07416_ (.A1(_01918_),
    .A2(_01921_),
    .B1(_01917_),
    .Y(_01970_));
 sky130_fd_sc_hd__xor2_4 _07417_ (.A(_01969_),
    .B(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__a221oi_1 _07418_ (.A1(_01965_),
    .A2(_01966_),
    .B1(_01971_),
    .B2(_01856_),
    .C1(_01884_),
    .Y(_01972_));
 sky130_fd_sc_hd__a211o_1 _07419_ (.A1(_01632_),
    .A2(_01827_),
    .B1(_01693_),
    .C1(_01972_),
    .X(_00252_));
 sky130_fd_sc_hd__buf_4 _07420_ (.A(_01421_),
    .X(_01973_));
 sky130_fd_sc_hd__inv_2 _07421_ (.A(_01952_),
    .Y(_01974_));
 sky130_fd_sc_hd__or2_1 _07422_ (.A(_01974_),
    .B(_01955_),
    .X(_01975_));
 sky130_fd_sc_hd__xnor2_1 _07423_ (.A(_01657_),
    .B(_01612_),
    .Y(_01976_));
 sky130_fd_sc_hd__xnor2_2 _07424_ (.A(_01675_),
    .B(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__or2_1 _07425_ (.A(\_185_[10] ),
    .B(\_234_[10] ),
    .X(_01978_));
 sky130_fd_sc_hd__nand2_1 _07426_ (.A(\_185_[10] ),
    .B(\_234_[10] ),
    .Y(_01979_));
 sky130_fd_sc_hd__nand2_1 _07427_ (.A(_01978_),
    .B(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__xor2_1 _07428_ (.A(_01977_),
    .B(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__a21o_1 _07429_ (.A1(_01954_),
    .A2(_01975_),
    .B1(_01981_),
    .X(_01982_));
 sky130_fd_sc_hd__nand3_1 _07430_ (.A(_01954_),
    .B(_01975_),
    .C(_01981_),
    .Y(_01983_));
 sky130_fd_sc_hd__nand2_1 _07431_ (.A(_01982_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__mux2_2 _07432_ (.A0(\_243_[10] ),
    .A1(\_240_[10] ),
    .S(_01635_),
    .X(_01985_));
 sky130_fd_sc_hd__xnor2_1 _07433_ (.A(_01984_),
    .B(_01985_),
    .Y(_01986_));
 sky130_fd_sc_hd__and2b_1 _07434_ (.A_N(_01959_),
    .B(_01960_),
    .X(_01987_));
 sky130_fd_sc_hd__or2_1 _07435_ (.A(_01957_),
    .B(_01987_),
    .X(_01988_));
 sky130_fd_sc_hd__nand2_1 _07436_ (.A(_01986_),
    .B(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__or2_1 _07437_ (.A(_01986_),
    .B(_01988_),
    .X(_01990_));
 sky130_fd_sc_hd__nand2_1 _07438_ (.A(_01989_),
    .B(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__or2b_1 _07439_ (.A(_01941_),
    .B_N(_01963_),
    .X(_01992_));
 sky130_fd_sc_hd__o21ai_1 _07440_ (.A1(_01944_),
    .A2(_01992_),
    .B1(_01962_),
    .Y(_01993_));
 sky130_fd_sc_hd__or2_1 _07441_ (.A(_01991_),
    .B(_01993_),
    .X(_01994_));
 sky130_fd_sc_hd__a21oi_1 _07442_ (.A1(_01991_),
    .A2(_01993_),
    .B1(_01409_),
    .Y(_01995_));
 sky130_fd_sc_hd__nand2_1 _07443_ (.A(\_182_[10] ),
    .B(_01635_),
    .Y(_01996_));
 sky130_fd_sc_hd__or2_1 _07444_ (.A(\_182_[10] ),
    .B(_01635_),
    .X(_01997_));
 sky130_fd_sc_hd__nand2_1 _07445_ (.A(_01996_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__nand3_1 _07446_ (.A(\_182_[8] ),
    .B(_01629_),
    .C(_01967_),
    .Y(_01999_));
 sky130_fd_sc_hd__o311a_1 _07447_ (.A1(_01918_),
    .A2(_01921_),
    .A3(_01969_),
    .B1(_01999_),
    .C1(_01968_),
    .X(_02000_));
 sky130_fd_sc_hd__xor2_2 _07448_ (.A(_01998_),
    .B(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__clkbuf_4 _07449_ (.A(_01404_),
    .X(_02002_));
 sky130_fd_sc_hd__a21o_1 _07450_ (.A1(_01923_),
    .A2(_02001_),
    .B1(_02002_),
    .X(_02003_));
 sky130_fd_sc_hd__a21o_1 _07451_ (.A1(_01994_),
    .A2(_01995_),
    .B1(_02003_),
    .X(_02004_));
 sky130_fd_sc_hd__o211a_1 _07452_ (.A1(_01635_),
    .A2(_01973_),
    .B1(_01886_),
    .C1(_02004_),
    .X(_00253_));
 sky130_fd_sc_hd__or2b_1 _07453_ (.A(_01984_),
    .B_N(_01985_),
    .X(_02005_));
 sky130_fd_sc_hd__inv_2 _07454_ (.A(_01977_),
    .Y(_02006_));
 sky130_fd_sc_hd__or2_1 _07455_ (.A(_02006_),
    .B(_01980_),
    .X(_02007_));
 sky130_fd_sc_hd__xnor2_1 _07456_ (.A(_01661_),
    .B(_01616_),
    .Y(_02008_));
 sky130_fd_sc_hd__xnor2_1 _07457_ (.A(_01678_),
    .B(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__or2_1 _07458_ (.A(\_185_[11] ),
    .B(\_234_[11] ),
    .X(_02010_));
 sky130_fd_sc_hd__nand2_1 _07459_ (.A(\_185_[11] ),
    .B(\_234_[11] ),
    .Y(_02011_));
 sky130_fd_sc_hd__nand2_1 _07460_ (.A(_02010_),
    .B(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hd__xor2_1 _07461_ (.A(_02009_),
    .B(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__a21oi_1 _07462_ (.A1(_01979_),
    .A2(_02007_),
    .B1(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__and3_1 _07463_ (.A(_01979_),
    .B(_02007_),
    .C(_02013_),
    .X(_02015_));
 sky130_fd_sc_hd__or2_1 _07464_ (.A(_02014_),
    .B(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_2 _07465_ (.A0(\_243_[11] ),
    .A1(\_240_[11] ),
    .S(_01638_),
    .X(_02017_));
 sky130_fd_sc_hd__xor2_1 _07466_ (.A(_02016_),
    .B(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__a21oi_1 _07467_ (.A1(_01982_),
    .A2(_02005_),
    .B1(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__nand3_1 _07468_ (.A(_01982_),
    .B(_02005_),
    .C(_02018_),
    .Y(_02020_));
 sky130_fd_sc_hd__or2b_1 _07469_ (.A(_02019_),
    .B_N(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__a21oi_1 _07470_ (.A1(_01989_),
    .A2(_01994_),
    .B1(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__a31o_1 _07471_ (.A1(_01989_),
    .A2(_01994_),
    .A3(_02021_),
    .B1(_01923_),
    .X(_02023_));
 sky130_fd_sc_hd__nand2_1 _07472_ (.A(\_182_[11] ),
    .B(_01638_),
    .Y(_02024_));
 sky130_fd_sc_hd__or2_1 _07473_ (.A(\_182_[11] ),
    .B(_01638_),
    .X(_02025_));
 sky130_fd_sc_hd__nand2_2 _07474_ (.A(_02024_),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__o21a_2 _07475_ (.A1(_01998_),
    .A2(_02000_),
    .B1(_01996_),
    .X(_02027_));
 sky130_fd_sc_hd__xor2_4 _07476_ (.A(_02026_),
    .B(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__a21oi_1 _07477_ (.A1(_01428_),
    .A2(_02028_),
    .B1(_01495_),
    .Y(_02029_));
 sky130_fd_sc_hd__o21ai_1 _07478_ (.A1(_02022_),
    .A2(_02023_),
    .B1(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__o211a_1 _07479_ (.A1(_01638_),
    .A2(_01973_),
    .B1(_01886_),
    .C1(_02030_),
    .X(_00254_));
 sky130_fd_sc_hd__nor2_1 _07480_ (.A(_01991_),
    .B(_02021_),
    .Y(_02031_));
 sky130_fd_sc_hd__o2111ai_4 _07481_ (.A1(_01924_),
    .A2(_01925_),
    .B1(_01964_),
    .C1(_02031_),
    .D1(_01943_),
    .Y(_02032_));
 sky130_fd_sc_hd__a31o_1 _07482_ (.A1(_01986_),
    .A2(_01988_),
    .A3(_02020_),
    .B1(_02019_),
    .X(_02033_));
 sky130_fd_sc_hd__a31oi_2 _07483_ (.A1(_01962_),
    .A2(_01992_),
    .A3(_02031_),
    .B1(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _07484_ (.A(_02032_),
    .B(_02034_),
    .Y(_02035_));
 sky130_fd_sc_hd__and2b_1 _07485_ (.A_N(_02016_),
    .B(_02017_),
    .X(_02036_));
 sky130_fd_sc_hd__inv_2 _07486_ (.A(_02009_),
    .Y(_02037_));
 sky130_fd_sc_hd__or2_1 _07487_ (.A(_02037_),
    .B(_02012_),
    .X(_02038_));
 sky130_fd_sc_hd__xnor2_1 _07488_ (.A(_01664_),
    .B(_01620_),
    .Y(_02039_));
 sky130_fd_sc_hd__xnor2_1 _07489_ (.A(_01681_),
    .B(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__or2_1 _07490_ (.A(\_185_[12] ),
    .B(\_234_[12] ),
    .X(_02041_));
 sky130_fd_sc_hd__nand2_1 _07491_ (.A(\_185_[12] ),
    .B(\_234_[12] ),
    .Y(_02042_));
 sky130_fd_sc_hd__nand2_1 _07492_ (.A(_02041_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__xor2_1 _07493_ (.A(_02040_),
    .B(_02043_),
    .X(_02044_));
 sky130_fd_sc_hd__a21oi_1 _07494_ (.A1(_02011_),
    .A2(_02038_),
    .B1(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__and3_1 _07495_ (.A(_02011_),
    .B(_02038_),
    .C(_02044_),
    .X(_02046_));
 sky130_fd_sc_hd__or2_1 _07496_ (.A(_02045_),
    .B(_02046_),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_2 _07497_ (.A0(\_243_[12] ),
    .A1(\_240_[12] ),
    .S(_01642_),
    .X(_02048_));
 sky130_fd_sc_hd__xnor2_1 _07498_ (.A(_02047_),
    .B(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__o21a_1 _07499_ (.A1(_02014_),
    .A2(_02036_),
    .B1(_02049_),
    .X(_02050_));
 sky130_fd_sc_hd__nor3_1 _07500_ (.A(_02014_),
    .B(_02036_),
    .C(_02049_),
    .Y(_02051_));
 sky130_fd_sc_hd__nor2_1 _07501_ (.A(_02050_),
    .B(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__xnor2_1 _07502_ (.A(_02035_),
    .B(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__o21a_1 _07503_ (.A1(_02026_),
    .A2(_02027_),
    .B1(_02024_),
    .X(_02054_));
 sky130_fd_sc_hd__xor2_1 _07504_ (.A(\_182_[12] ),
    .B(_01642_),
    .X(_02055_));
 sky130_fd_sc_hd__and2b_1 _07505_ (.A_N(_02054_),
    .B(_02055_),
    .X(_02056_));
 sky130_fd_sc_hd__and2b_1 _07506_ (.A_N(_02055_),
    .B(_02054_),
    .X(_02057_));
 sky130_fd_sc_hd__or2_2 _07507_ (.A(_02056_),
    .B(_02057_),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _07508_ (.A0(_02053_),
    .A1(_02058_),
    .S(_01427_),
    .X(_02059_));
 sky130_fd_sc_hd__nor2_1 _07509_ (.A(_01884_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__a211o_1 _07510_ (.A1(_01642_),
    .A2(_01827_),
    .B1(_01693_),
    .C1(_02060_),
    .X(_00255_));
 sky130_fd_sc_hd__and2b_1 _07511_ (.A_N(_02047_),
    .B(_02048_),
    .X(_02061_));
 sky130_fd_sc_hd__xnor2_1 _07512_ (.A(_01667_),
    .B(_01623_),
    .Y(_02062_));
 sky130_fd_sc_hd__xnor2_1 _07513_ (.A(_01684_),
    .B(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__inv_2 _07514_ (.A(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__or2_1 _07515_ (.A(\_185_[13] ),
    .B(\_234_[13] ),
    .X(_02065_));
 sky130_fd_sc_hd__nand2_1 _07516_ (.A(\_185_[13] ),
    .B(\_234_[13] ),
    .Y(_02066_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(_02065_),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__or2_1 _07518_ (.A(_02064_),
    .B(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__nand2_1 _07519_ (.A(_02064_),
    .B(_02067_),
    .Y(_02069_));
 sky130_fd_sc_hd__nand2_1 _07520_ (.A(_02068_),
    .B(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__inv_2 _07521_ (.A(_02040_),
    .Y(_02071_));
 sky130_fd_sc_hd__o21a_1 _07522_ (.A1(_02071_),
    .A2(_02043_),
    .B1(_02042_),
    .X(_02072_));
 sky130_fd_sc_hd__xnor2_1 _07523_ (.A(_02070_),
    .B(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__mux2_2 _07524_ (.A0(\_243_[13] ),
    .A1(\_240_[13] ),
    .S(_01645_),
    .X(_02074_));
 sky130_fd_sc_hd__xnor2_1 _07525_ (.A(_02073_),
    .B(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__o21a_1 _07526_ (.A1(_02045_),
    .A2(_02061_),
    .B1(_02075_),
    .X(_02076_));
 sky130_fd_sc_hd__or3_2 _07527_ (.A(_02045_),
    .B(_02061_),
    .C(_02075_),
    .X(_02077_));
 sky130_fd_sc_hd__and2b_1 _07528_ (.A_N(_02076_),
    .B(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__a21oi_1 _07529_ (.A1(_02035_),
    .A2(_02052_),
    .B1(_02050_),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_1 _07530_ (.A(_02078_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__or2_1 _07531_ (.A(\_182_[13] ),
    .B(_01645_),
    .X(_02081_));
 sky130_fd_sc_hd__nand2_1 _07532_ (.A(\_182_[13] ),
    .B(_01645_),
    .Y(_02082_));
 sky130_fd_sc_hd__nand2_1 _07533_ (.A(_02081_),
    .B(_02082_),
    .Y(_02083_));
 sky130_fd_sc_hd__a21oi_1 _07534_ (.A1(\_182_[12] ),
    .A2(_01642_),
    .B1(_02056_),
    .Y(_02084_));
 sky130_fd_sc_hd__xnor2_2 _07535_ (.A(_02083_),
    .B(_02084_),
    .Y(_02085_));
 sky130_fd_sc_hd__nor2_1 _07536_ (.A(_01778_),
    .B(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__a211o_1 _07537_ (.A1(_01355_),
    .A2(_02080_),
    .B1(_02086_),
    .C1(_01884_),
    .X(_02087_));
 sky130_fd_sc_hd__o211a_1 _07538_ (.A1(_01645_),
    .A2(_01973_),
    .B1(_01886_),
    .C1(_02087_),
    .X(_00256_));
 sky130_fd_sc_hd__xnor2_1 _07539_ (.A(_01671_),
    .B(_01626_),
    .Y(_02088_));
 sky130_fd_sc_hd__xnor2_1 _07540_ (.A(_01687_),
    .B(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__or2_1 _07541_ (.A(\_185_[14] ),
    .B(\_234_[14] ),
    .X(_02090_));
 sky130_fd_sc_hd__nand2_1 _07542_ (.A(\_185_[14] ),
    .B(\_234_[14] ),
    .Y(_02091_));
 sky130_fd_sc_hd__nand2_1 _07543_ (.A(_02090_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__xor2_1 _07544_ (.A(_02089_),
    .B(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__a21oi_1 _07545_ (.A1(_02066_),
    .A2(_02068_),
    .B1(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__and3_1 _07546_ (.A(_02066_),
    .B(_02068_),
    .C(_02093_),
    .X(_02095_));
 sky130_fd_sc_hd__or2_1 _07547_ (.A(_02094_),
    .B(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__mux2_2 _07548_ (.A0(\_243_[14] ),
    .A1(\_240_[14] ),
    .S(_01650_),
    .X(_02097_));
 sky130_fd_sc_hd__xnor2_1 _07549_ (.A(_02096_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__and2b_1 _07550_ (.A_N(_02073_),
    .B(_02074_),
    .X(_02099_));
 sky130_fd_sc_hd__o21ba_1 _07551_ (.A1(_02070_),
    .A2(_02072_),
    .B1_N(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__xnor2_1 _07552_ (.A(_02098_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__or2_1 _07553_ (.A(_02050_),
    .B(_02076_),
    .X(_02102_));
 sky130_fd_sc_hd__and2_1 _07554_ (.A(_02077_),
    .B(_02102_),
    .X(_02103_));
 sky130_fd_sc_hd__a31o_1 _07555_ (.A1(_02035_),
    .A2(_02052_),
    .A3(_02078_),
    .B1(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__xor2_1 _07556_ (.A(_02101_),
    .B(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__or2_1 _07557_ (.A(\_182_[14] ),
    .B(_01650_),
    .X(_02106_));
 sky130_fd_sc_hd__nand2_1 _07558_ (.A(\_182_[14] ),
    .B(_01650_),
    .Y(_02107_));
 sky130_fd_sc_hd__nand2_1 _07559_ (.A(_02106_),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__a22o_1 _07560_ (.A1(\_182_[13] ),
    .A2(_01645_),
    .B1(_01642_),
    .B2(\_182_[12] ),
    .X(_02109_));
 sky130_fd_sc_hd__o21ai_2 _07561_ (.A1(_02056_),
    .A2(_02109_),
    .B1(_02081_),
    .Y(_02110_));
 sky130_fd_sc_hd__xnor2_2 _07562_ (.A(_02108_),
    .B(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__nand2_1 _07563_ (.A(_01409_),
    .B(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__o211a_1 _07564_ (.A1(_01801_),
    .A2(_02105_),
    .B1(_02112_),
    .C1(_01799_),
    .X(_02113_));
 sky130_fd_sc_hd__a211o_1 _07565_ (.A1(_01650_),
    .A2(_01827_),
    .B1(_01693_),
    .C1(_02113_),
    .X(_00257_));
 sky130_fd_sc_hd__and2b_1 _07566_ (.A_N(_02096_),
    .B(_02097_),
    .X(_02114_));
 sky130_fd_sc_hd__xnor2_1 _07567_ (.A(_01675_),
    .B(_01629_),
    .Y(_02115_));
 sky130_fd_sc_hd__xnor2_1 _07568_ (.A(_01690_),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__inv_2 _07569_ (.A(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__or2_1 _07570_ (.A(\_185_[15] ),
    .B(\_234_[15] ),
    .X(_02118_));
 sky130_fd_sc_hd__nand2_1 _07571_ (.A(\_185_[15] ),
    .B(\_234_[15] ),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_1 _07572_ (.A(_02118_),
    .B(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__or2_1 _07573_ (.A(_02117_),
    .B(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__nand2_1 _07574_ (.A(_02117_),
    .B(_02120_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_1 _07575_ (.A(_02121_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__inv_2 _07576_ (.A(_02089_),
    .Y(_02124_));
 sky130_fd_sc_hd__o21a_1 _07577_ (.A1(_02124_),
    .A2(_02092_),
    .B1(_02091_),
    .X(_02125_));
 sky130_fd_sc_hd__xnor2_1 _07578_ (.A(_02123_),
    .B(_02125_),
    .Y(_02126_));
 sky130_fd_sc_hd__mux2_4 _07579_ (.A0(\_243_[15] ),
    .A1(\_240_[15] ),
    .S(_01654_),
    .X(_02127_));
 sky130_fd_sc_hd__xnor2_1 _07580_ (.A(_02126_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__o21a_1 _07581_ (.A1(_02094_),
    .A2(_02114_),
    .B1(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__nor3_1 _07582_ (.A(_02094_),
    .B(_02114_),
    .C(_02128_),
    .Y(_02130_));
 sky130_fd_sc_hd__nor2_1 _07583_ (.A(_02129_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__or2b_1 _07584_ (.A(_02100_),
    .B_N(_02098_),
    .X(_02132_));
 sky130_fd_sc_hd__a21bo_1 _07585_ (.A1(_02101_),
    .A2(_02104_),
    .B1_N(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__xnor2_1 _07586_ (.A(_02131_),
    .B(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__nor2_1 _07587_ (.A(\_182_[15] ),
    .B(_01654_),
    .Y(_02135_));
 sky130_fd_sc_hd__nand2_1 _07588_ (.A(\_182_[15] ),
    .B(_01654_),
    .Y(_02136_));
 sky130_fd_sc_hd__and2b_1 _07589_ (.A_N(_02135_),
    .B(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__o21ai_1 _07590_ (.A1(_02108_),
    .A2(_02110_),
    .B1(_02107_),
    .Y(_02138_));
 sky130_fd_sc_hd__xnor2_2 _07591_ (.A(_02137_),
    .B(_02138_),
    .Y(_02139_));
 sky130_fd_sc_hd__mux2_1 _07592_ (.A0(_02134_),
    .A1(_02139_),
    .S(_01427_),
    .X(_02140_));
 sky130_fd_sc_hd__nand2_1 _07593_ (.A(_01444_),
    .B(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__o211a_1 _07594_ (.A1(_01654_),
    .A2(_01973_),
    .B1(_01886_),
    .C1(_02141_),
    .X(_00258_));
 sky130_fd_sc_hd__and2_1 _07595_ (.A(_02101_),
    .B(_02131_),
    .X(_02142_));
 sky130_fd_sc_hd__nor2_1 _07596_ (.A(_02132_),
    .B(_02130_),
    .Y(_02143_));
 sky130_fd_sc_hd__a311oi_4 _07597_ (.A1(_02077_),
    .A2(_02102_),
    .A3(_02142_),
    .B1(_02143_),
    .C1(_02129_),
    .Y(_02144_));
 sky130_fd_sc_hd__nand2_1 _07598_ (.A(_02052_),
    .B(_02078_),
    .Y(_02145_));
 sky130_fd_sc_hd__inv_2 _07599_ (.A(_02142_),
    .Y(_02146_));
 sky130_fd_sc_hd__a211o_1 _07600_ (.A1(_02032_),
    .A2(_02034_),
    .B1(_02145_),
    .C1(_02146_),
    .X(_02147_));
 sky130_fd_sc_hd__nand2_1 _07601_ (.A(_02144_),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__xnor2_1 _07602_ (.A(_01678_),
    .B(_01632_),
    .Y(_02149_));
 sky130_fd_sc_hd__xnor2_1 _07603_ (.A(_01694_),
    .B(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__inv_2 _07604_ (.A(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__or2_1 _07605_ (.A(\_185_[16] ),
    .B(\_234_[16] ),
    .X(_02152_));
 sky130_fd_sc_hd__nand2_1 _07606_ (.A(\_185_[16] ),
    .B(\_234_[16] ),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2_1 _07607_ (.A(_02152_),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__or2_1 _07608_ (.A(_02151_),
    .B(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__nand2_1 _07609_ (.A(_02151_),
    .B(_02154_),
    .Y(_02156_));
 sky130_fd_sc_hd__nand2_1 _07610_ (.A(_02155_),
    .B(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__a21oi_1 _07611_ (.A1(_02119_),
    .A2(_02121_),
    .B1(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__and3_1 _07612_ (.A(_02119_),
    .B(_02121_),
    .C(_02157_),
    .X(_02159_));
 sky130_fd_sc_hd__or2_1 _07613_ (.A(_02158_),
    .B(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__mux2_4 _07614_ (.A0(\_243_[16] ),
    .A1(\_240_[16] ),
    .S(_01657_),
    .X(_02161_));
 sky130_fd_sc_hd__xnor2_1 _07615_ (.A(_02160_),
    .B(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__and2b_1 _07616_ (.A_N(_02126_),
    .B(_02127_),
    .X(_02163_));
 sky130_fd_sc_hd__o21ba_1 _07617_ (.A1(_02123_),
    .A2(_02125_),
    .B1_N(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__xnor2_1 _07618_ (.A(_02162_),
    .B(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__nand2_1 _07619_ (.A(_02148_),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__or2_1 _07620_ (.A(_02148_),
    .B(_02165_),
    .X(_02167_));
 sky130_fd_sc_hd__nor2_1 _07621_ (.A(\_182_[16] ),
    .B(_01657_),
    .Y(_02168_));
 sky130_fd_sc_hd__and2_1 _07622_ (.A(\_182_[16] ),
    .B(_01657_),
    .X(_02169_));
 sky130_fd_sc_hd__or2_1 _07623_ (.A(_02168_),
    .B(_02169_),
    .X(_02170_));
 sky130_fd_sc_hd__nand3b_1 _07624_ (.A_N(_02135_),
    .B(_01650_),
    .C(\_182_[14] ),
    .Y(_02171_));
 sky130_fd_sc_hd__o311a_1 _07625_ (.A1(_02108_),
    .A2(_02110_),
    .A3(_02135_),
    .B1(_02136_),
    .C1(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__nor2_1 _07626_ (.A(_02170_),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__and2_1 _07627_ (.A(_02170_),
    .B(_02172_),
    .X(_02174_));
 sky130_fd_sc_hd__nor2_2 _07628_ (.A(_02173_),
    .B(_02174_),
    .Y(_02175_));
 sky130_fd_sc_hd__a21o_1 _07629_ (.A1(_01923_),
    .A2(_02175_),
    .B1(_02002_),
    .X(_02176_));
 sky130_fd_sc_hd__a31o_1 _07630_ (.A1(_01355_),
    .A2(_02166_),
    .A3(_02167_),
    .B1(_02176_),
    .X(_02177_));
 sky130_fd_sc_hd__o211a_1 _07631_ (.A1(_01657_),
    .A2(_01973_),
    .B1(_01886_),
    .C1(_02177_),
    .X(_00259_));
 sky130_fd_sc_hd__buf_2 _07632_ (.A(_01435_),
    .X(_02178_));
 sky130_fd_sc_hd__xnor2_2 _07633_ (.A(\_182_[17] ),
    .B(_01661_),
    .Y(_02179_));
 sky130_fd_sc_hd__or2_2 _07634_ (.A(_02169_),
    .B(_02173_),
    .X(_02180_));
 sky130_fd_sc_hd__xnor2_4 _07635_ (.A(_02179_),
    .B(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__and2b_1 _07636_ (.A_N(_02160_),
    .B(_02161_),
    .X(_02182_));
 sky130_fd_sc_hd__xnor2_1 _07637_ (.A(_01681_),
    .B(_01635_),
    .Y(_02183_));
 sky130_fd_sc_hd__xnor2_2 _07638_ (.A(_01698_),
    .B(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__or2_1 _07639_ (.A(\_185_[17] ),
    .B(\_234_[17] ),
    .X(_02185_));
 sky130_fd_sc_hd__nand2_1 _07640_ (.A(\_185_[17] ),
    .B(\_234_[17] ),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_1 _07641_ (.A(_02185_),
    .B(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__xor2_1 _07642_ (.A(_02184_),
    .B(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__a21oi_1 _07643_ (.A1(_02153_),
    .A2(_02155_),
    .B1(_02188_),
    .Y(_02189_));
 sky130_fd_sc_hd__and3_1 _07644_ (.A(_02153_),
    .B(_02155_),
    .C(_02188_),
    .X(_02190_));
 sky130_fd_sc_hd__or2_1 _07645_ (.A(_02189_),
    .B(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_4 _07646_ (.A0(\_243_[17] ),
    .A1(\_240_[17] ),
    .S(_01661_),
    .X(_02192_));
 sky130_fd_sc_hd__xnor2_1 _07647_ (.A(_02191_),
    .B(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__o21ai_1 _07648_ (.A1(_02158_),
    .A2(_02182_),
    .B1(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__inv_2 _07649_ (.A(_02194_),
    .Y(_02195_));
 sky130_fd_sc_hd__nor3_1 _07650_ (.A(_02158_),
    .B(_02182_),
    .C(_02193_),
    .Y(_02196_));
 sky130_fd_sc_hd__nor2_1 _07651_ (.A(_02195_),
    .B(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__or2b_1 _07652_ (.A(_02164_),
    .B_N(_02162_),
    .X(_02198_));
 sky130_fd_sc_hd__and2_1 _07653_ (.A(_02198_),
    .B(_02166_),
    .X(_02199_));
 sky130_fd_sc_hd__o21ai_1 _07654_ (.A1(_02197_),
    .A2(_02199_),
    .B1(_01519_),
    .Y(_02200_));
 sky130_fd_sc_hd__a21o_1 _07655_ (.A1(_02197_),
    .A2(_02199_),
    .B1(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__clkbuf_4 _07656_ (.A(_01412_),
    .X(_02202_));
 sky130_fd_sc_hd__o211a_1 _07657_ (.A1(_01520_),
    .A2(_02181_),
    .B1(_02201_),
    .C1(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__a211o_1 _07658_ (.A1(_01661_),
    .A2(_01827_),
    .B1(_02178_),
    .C1(_02203_),
    .X(_00260_));
 sky130_fd_sc_hd__and2b_1 _07659_ (.A_N(_02191_),
    .B(_02192_),
    .X(_02204_));
 sky130_fd_sc_hd__inv_2 _07660_ (.A(_02184_),
    .Y(_02205_));
 sky130_fd_sc_hd__or2_1 _07661_ (.A(_02205_),
    .B(_02187_),
    .X(_02206_));
 sky130_fd_sc_hd__xnor2_2 _07662_ (.A(_01684_),
    .B(_01638_),
    .Y(_02207_));
 sky130_fd_sc_hd__xnor2_2 _07663_ (.A(_01701_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__or2_1 _07664_ (.A(\_185_[18] ),
    .B(\_234_[18] ),
    .X(_02209_));
 sky130_fd_sc_hd__nand2_1 _07665_ (.A(\_185_[18] ),
    .B(\_234_[18] ),
    .Y(_02210_));
 sky130_fd_sc_hd__nand2_1 _07666_ (.A(_02209_),
    .B(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__xor2_1 _07667_ (.A(_02208_),
    .B(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__a21oi_1 _07668_ (.A1(_02186_),
    .A2(_02206_),
    .B1(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__and3_1 _07669_ (.A(_02186_),
    .B(_02206_),
    .C(_02212_),
    .X(_02214_));
 sky130_fd_sc_hd__or2_1 _07670_ (.A(_02213_),
    .B(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__mux2_4 _07671_ (.A0(\_243_[18] ),
    .A1(\_240_[18] ),
    .S(_01664_),
    .X(_02216_));
 sky130_fd_sc_hd__xnor2_1 _07672_ (.A(_02215_),
    .B(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__o21ai_1 _07673_ (.A1(_02189_),
    .A2(_02204_),
    .B1(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__or3_1 _07674_ (.A(_02189_),
    .B(_02204_),
    .C(_02217_),
    .X(_02219_));
 sky130_fd_sc_hd__and2_1 _07675_ (.A(_02218_),
    .B(_02219_),
    .X(_02220_));
 sky130_fd_sc_hd__inv_2 _07676_ (.A(_02197_),
    .Y(_02221_));
 sky130_fd_sc_hd__a21o_1 _07677_ (.A1(_02198_),
    .A2(_02194_),
    .B1(_02196_),
    .X(_02222_));
 sky130_fd_sc_hd__o21ai_2 _07678_ (.A1(_02166_),
    .A2(_02221_),
    .B1(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__xor2_2 _07679_ (.A(_02220_),
    .B(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__nor2_1 _07680_ (.A(\_182_[18] ),
    .B(_01664_),
    .Y(_02225_));
 sky130_fd_sc_hd__and2_1 _07681_ (.A(\_182_[18] ),
    .B(_01664_),
    .X(_02226_));
 sky130_fd_sc_hd__nor2_2 _07682_ (.A(_02225_),
    .B(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__a21o_1 _07683_ (.A1(\_182_[17] ),
    .A2(_01661_),
    .B1(_02169_),
    .X(_02228_));
 sky130_fd_sc_hd__o22a_2 _07684_ (.A1(\_182_[17] ),
    .A2(_01661_),
    .B1(_02173_),
    .B2(_02228_),
    .X(_02229_));
 sky130_fd_sc_hd__xnor2_4 _07685_ (.A(_02227_),
    .B(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hd__nand2_1 _07686_ (.A(_01409_),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__o211a_1 _07687_ (.A1(_01801_),
    .A2(_02224_),
    .B1(_02231_),
    .C1(_02202_),
    .X(_02232_));
 sky130_fd_sc_hd__a211o_1 _07688_ (.A1(_01664_),
    .A2(_01827_),
    .B1(_02178_),
    .C1(_02232_),
    .X(_00261_));
 sky130_fd_sc_hd__nor2_1 _07689_ (.A(\_182_[19] ),
    .B(_01667_),
    .Y(_02233_));
 sky130_fd_sc_hd__nand2_1 _07690_ (.A(\_182_[19] ),
    .B(_01667_),
    .Y(_02234_));
 sky130_fd_sc_hd__and2b_2 _07691_ (.A_N(_02233_),
    .B(_02234_),
    .X(_02235_));
 sky130_fd_sc_hd__a21oi_2 _07692_ (.A1(_02227_),
    .A2(_02229_),
    .B1(_02226_),
    .Y(_02236_));
 sky130_fd_sc_hd__xnor2_4 _07693_ (.A(_02235_),
    .B(_02236_),
    .Y(_02237_));
 sky130_fd_sc_hd__nand2_1 _07694_ (.A(_02220_),
    .B(_02223_),
    .Y(_02238_));
 sky130_fd_sc_hd__and2b_1 _07695_ (.A_N(_02215_),
    .B(_02216_),
    .X(_02239_));
 sky130_fd_sc_hd__xnor2_1 _07696_ (.A(_01687_),
    .B(_01642_),
    .Y(_02240_));
 sky130_fd_sc_hd__xnor2_1 _07697_ (.A(_01704_),
    .B(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__inv_2 _07698_ (.A(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__or2_1 _07699_ (.A(\_185_[19] ),
    .B(\_234_[19] ),
    .X(_02243_));
 sky130_fd_sc_hd__nand2_1 _07700_ (.A(\_185_[19] ),
    .B(\_234_[19] ),
    .Y(_02244_));
 sky130_fd_sc_hd__nand2_1 _07701_ (.A(_02243_),
    .B(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__or2_1 _07702_ (.A(_02242_),
    .B(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__nand2_1 _07703_ (.A(_02242_),
    .B(_02245_),
    .Y(_02247_));
 sky130_fd_sc_hd__nand2_1 _07704_ (.A(_02246_),
    .B(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__inv_2 _07705_ (.A(_02208_),
    .Y(_02249_));
 sky130_fd_sc_hd__o21a_1 _07706_ (.A1(_02249_),
    .A2(_02211_),
    .B1(_02210_),
    .X(_02250_));
 sky130_fd_sc_hd__xnor2_1 _07707_ (.A(_02248_),
    .B(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__mux2_4 _07708_ (.A0(\_243_[19] ),
    .A1(\_240_[19] ),
    .S(_01667_),
    .X(_02252_));
 sky130_fd_sc_hd__xnor2_1 _07709_ (.A(_02251_),
    .B(_02252_),
    .Y(_02253_));
 sky130_fd_sc_hd__o21a_1 _07710_ (.A1(_02213_),
    .A2(_02239_),
    .B1(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__nor3_1 _07711_ (.A(_02213_),
    .B(_02239_),
    .C(_02253_),
    .Y(_02255_));
 sky130_fd_sc_hd__nor2_1 _07712_ (.A(_02254_),
    .B(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__a21oi_1 _07713_ (.A1(_02218_),
    .A2(_02238_),
    .B1(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__a31o_1 _07714_ (.A1(_02218_),
    .A2(_02238_),
    .A3(_02256_),
    .B1(_01269_),
    .X(_02258_));
 sky130_fd_sc_hd__or2_1 _07715_ (.A(_02257_),
    .B(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__o211a_1 _07716_ (.A1(_01520_),
    .A2(_02237_),
    .B1(_02259_),
    .C1(_02202_),
    .X(_02260_));
 sky130_fd_sc_hd__a211o_1 _07717_ (.A1(_01667_),
    .A2(_01827_),
    .B1(_02178_),
    .C1(_02260_),
    .X(_00262_));
 sky130_fd_sc_hd__xnor2_2 _07718_ (.A(_01690_),
    .B(_01645_),
    .Y(_02261_));
 sky130_fd_sc_hd__xnor2_4 _07719_ (.A(_01707_),
    .B(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__or2_1 _07720_ (.A(\_185_[20] ),
    .B(\_234_[20] ),
    .X(_02263_));
 sky130_fd_sc_hd__nand2_1 _07721_ (.A(\_185_[20] ),
    .B(\_234_[20] ),
    .Y(_02264_));
 sky130_fd_sc_hd__nand3_1 _07722_ (.A(_02262_),
    .B(_02263_),
    .C(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__a21o_1 _07723_ (.A1(_02263_),
    .A2(_02264_),
    .B1(_02262_),
    .X(_02266_));
 sky130_fd_sc_hd__nand2_1 _07724_ (.A(_02265_),
    .B(_02266_),
    .Y(_02267_));
 sky130_fd_sc_hd__a21oi_1 _07725_ (.A1(_02244_),
    .A2(_02246_),
    .B1(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__and3_1 _07726_ (.A(_02244_),
    .B(_02246_),
    .C(_02267_),
    .X(_02269_));
 sky130_fd_sc_hd__or2_1 _07727_ (.A(_02268_),
    .B(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_4 _07728_ (.A0(\_243_[20] ),
    .A1(\_240_[20] ),
    .S(_01671_),
    .X(_02271_));
 sky130_fd_sc_hd__xnor2_1 _07729_ (.A(_02270_),
    .B(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__and2b_1 _07730_ (.A_N(_02251_),
    .B(_02252_),
    .X(_02273_));
 sky130_fd_sc_hd__o21ba_1 _07731_ (.A1(_02248_),
    .A2(_02250_),
    .B1_N(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__xnor2_1 _07732_ (.A(_02272_),
    .B(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hd__nand2_1 _07733_ (.A(_02220_),
    .B(_02256_),
    .Y(_02276_));
 sky130_fd_sc_hd__or4b_1 _07734_ (.A(_02195_),
    .B(_02196_),
    .C(_02276_),
    .D_N(_02165_),
    .X(_02277_));
 sky130_fd_sc_hd__inv_2 _07735_ (.A(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__o22ai_1 _07736_ (.A1(_02218_),
    .A2(_02255_),
    .B1(_02276_),
    .B2(_02222_),
    .Y(_02279_));
 sky130_fd_sc_hd__nor2_1 _07737_ (.A(_02254_),
    .B(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__a21bo_1 _07738_ (.A1(_02148_),
    .A2(_02278_),
    .B1_N(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__xor2_1 _07739_ (.A(_02275_),
    .B(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__nand2_1 _07740_ (.A(\_182_[18] ),
    .B(_01664_),
    .Y(_02283_));
 sky130_fd_sc_hd__o2111ai_1 _07741_ (.A1(\_182_[17] ),
    .A2(_01661_),
    .B1(_02227_),
    .C1(_02228_),
    .D1(_02235_),
    .Y(_02284_));
 sky130_fd_sc_hd__o211a_1 _07742_ (.A1(_02283_),
    .A2(_02233_),
    .B1(_02234_),
    .C1(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__or4bb_1 _07743_ (.A(_02170_),
    .B(_02179_),
    .C_N(_02227_),
    .D_N(_02235_),
    .X(_02286_));
 sky130_fd_sc_hd__or2_1 _07744_ (.A(_02172_),
    .B(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__or2_1 _07745_ (.A(\_182_[20] ),
    .B(_01671_),
    .X(_02288_));
 sky130_fd_sc_hd__nand2_1 _07746_ (.A(\_182_[20] ),
    .B(_01671_),
    .Y(_02289_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(_02288_),
    .B(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__a21oi_1 _07748_ (.A1(_02285_),
    .A2(_02287_),
    .B1(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__and3_1 _07749_ (.A(_02290_),
    .B(_02285_),
    .C(_02287_),
    .X(_02292_));
 sky130_fd_sc_hd__or2_2 _07750_ (.A(_02291_),
    .B(_02292_),
    .X(_02293_));
 sky130_fd_sc_hd__nor2_1 _07751_ (.A(_01778_),
    .B(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__a211o_1 _07752_ (.A1(_01355_),
    .A2(_02282_),
    .B1(_02294_),
    .C1(_01884_),
    .X(_02295_));
 sky130_fd_sc_hd__o211a_1 _07753_ (.A1(_01671_),
    .A2(_01973_),
    .B1(_01886_),
    .C1(_02295_),
    .X(_00263_));
 sky130_fd_sc_hd__nand2_1 _07754_ (.A(\_182_[21] ),
    .B(_01675_),
    .Y(_02296_));
 sky130_fd_sc_hd__or2_1 _07755_ (.A(\_182_[21] ),
    .B(_01675_),
    .X(_02297_));
 sky130_fd_sc_hd__nand2_2 _07756_ (.A(_02296_),
    .B(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__a21o_1 _07757_ (.A1(\_182_[20] ),
    .A2(_01671_),
    .B1(_02291_),
    .X(_02299_));
 sky130_fd_sc_hd__xnor2_4 _07758_ (.A(_02298_),
    .B(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__and2b_1 _07759_ (.A_N(_02270_),
    .B(_02271_),
    .X(_02301_));
 sky130_fd_sc_hd__xnor2_2 _07760_ (.A(_01650_),
    .B(\_237_[0] ),
    .Y(_02302_));
 sky130_fd_sc_hd__xnor2_2 _07761_ (.A(_01694_),
    .B(_02302_),
    .Y(_02303_));
 sky130_fd_sc_hd__or2_1 _07762_ (.A(\_185_[21] ),
    .B(\_234_[21] ),
    .X(_02304_));
 sky130_fd_sc_hd__nand2_1 _07763_ (.A(\_185_[21] ),
    .B(\_234_[21] ),
    .Y(_02305_));
 sky130_fd_sc_hd__nand2_1 _07764_ (.A(_02304_),
    .B(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__xor2_1 _07765_ (.A(_02303_),
    .B(_02306_),
    .X(_02307_));
 sky130_fd_sc_hd__a21oi_1 _07766_ (.A1(_02264_),
    .A2(_02265_),
    .B1(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__and3_1 _07767_ (.A(_02264_),
    .B(_02265_),
    .C(_02307_),
    .X(_02309_));
 sky130_fd_sc_hd__or2_1 _07768_ (.A(_02308_),
    .B(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_4 _07769_ (.A0(\_243_[21] ),
    .A1(\_240_[21] ),
    .S(_01675_),
    .X(_02311_));
 sky130_fd_sc_hd__xnor2_1 _07770_ (.A(_02310_),
    .B(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__o21ai_1 _07771_ (.A1(_02268_),
    .A2(_02301_),
    .B1(_02312_),
    .Y(_02313_));
 sky130_fd_sc_hd__inv_2 _07772_ (.A(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__nor3_1 _07773_ (.A(_02268_),
    .B(_02301_),
    .C(_02312_),
    .Y(_02315_));
 sky130_fd_sc_hd__nor2_1 _07774_ (.A(_02314_),
    .B(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__or2b_1 _07775_ (.A(_02274_),
    .B_N(_02272_),
    .X(_02317_));
 sky130_fd_sc_hd__a21bo_1 _07776_ (.A1(_02275_),
    .A2(_02281_),
    .B1_N(_02317_),
    .X(_02318_));
 sky130_fd_sc_hd__a21oi_1 _07777_ (.A1(_02316_),
    .A2(_02318_),
    .B1(_01408_),
    .Y(_02319_));
 sky130_fd_sc_hd__o21a_1 _07778_ (.A1(_02316_),
    .A2(_02318_),
    .B1(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__a211o_1 _07779_ (.A1(_01856_),
    .A2(_02300_),
    .B1(_02320_),
    .C1(_01884_),
    .X(_02321_));
 sky130_fd_sc_hd__o211a_1 _07780_ (.A1(_01675_),
    .A2(_01973_),
    .B1(_01886_),
    .C1(_02321_),
    .X(_00264_));
 sky130_fd_sc_hd__and2b_1 _07781_ (.A_N(_02310_),
    .B(_02311_),
    .X(_02322_));
 sky130_fd_sc_hd__inv_2 _07782_ (.A(_02303_),
    .Y(_02323_));
 sky130_fd_sc_hd__or2_1 _07783_ (.A(_02323_),
    .B(_02306_),
    .X(_02324_));
 sky130_fd_sc_hd__xnor2_1 _07784_ (.A(_01654_),
    .B(_01604_),
    .Y(_02325_));
 sky130_fd_sc_hd__xnor2_2 _07785_ (.A(_01698_),
    .B(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__inv_2 _07786_ (.A(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__or2_1 _07787_ (.A(\_185_[22] ),
    .B(\_234_[22] ),
    .X(_02328_));
 sky130_fd_sc_hd__nand2_1 _07788_ (.A(\_185_[22] ),
    .B(\_234_[22] ),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_1 _07789_ (.A(_02328_),
    .B(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__or2_1 _07790_ (.A(_02327_),
    .B(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__nand2_1 _07791_ (.A(_02327_),
    .B(_02330_),
    .Y(_02332_));
 sky130_fd_sc_hd__nand2_1 _07792_ (.A(_02331_),
    .B(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__a21oi_1 _07793_ (.A1(_02305_),
    .A2(_02324_),
    .B1(_02333_),
    .Y(_02334_));
 sky130_fd_sc_hd__and3_1 _07794_ (.A(_02305_),
    .B(_02324_),
    .C(_02333_),
    .X(_02335_));
 sky130_fd_sc_hd__or2_1 _07795_ (.A(_02334_),
    .B(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__mux2_4 _07796_ (.A0(\_243_[22] ),
    .A1(\_240_[22] ),
    .S(_01678_),
    .X(_02337_));
 sky130_fd_sc_hd__xnor2_1 _07797_ (.A(_02336_),
    .B(_02337_),
    .Y(_02338_));
 sky130_fd_sc_hd__o21ai_1 _07798_ (.A1(_02308_),
    .A2(_02322_),
    .B1(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__or3_1 _07799_ (.A(_02308_),
    .B(_02322_),
    .C(_02338_),
    .X(_02340_));
 sky130_fd_sc_hd__and2_1 _07800_ (.A(_02339_),
    .B(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__nand2_1 _07801_ (.A(_02275_),
    .B(_02316_),
    .Y(_02342_));
 sky130_fd_sc_hd__inv_2 _07802_ (.A(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__a21o_1 _07803_ (.A1(_02317_),
    .A2(_02313_),
    .B1(_02315_),
    .X(_02344_));
 sky130_fd_sc_hd__a21bo_1 _07804_ (.A1(_02281_),
    .A2(_02343_),
    .B1_N(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__nand2_1 _07805_ (.A(_02341_),
    .B(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__o21a_1 _07806_ (.A1(_02341_),
    .A2(_02345_),
    .B1(_01354_),
    .X(_02347_));
 sky130_fd_sc_hd__nor2_1 _07807_ (.A(\_182_[22] ),
    .B(_01678_),
    .Y(_02348_));
 sky130_fd_sc_hd__and2_1 _07808_ (.A(\_182_[22] ),
    .B(_01678_),
    .X(_02349_));
 sky130_fd_sc_hd__nor2_2 _07809_ (.A(_02348_),
    .B(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__nand2_1 _07810_ (.A(_02289_),
    .B(_02296_),
    .Y(_02351_));
 sky130_fd_sc_hd__o21a_1 _07811_ (.A1(_02291_),
    .A2(_02351_),
    .B1(_02297_),
    .X(_02352_));
 sky130_fd_sc_hd__xor2_2 _07812_ (.A(_02350_),
    .B(_02352_),
    .X(_02353_));
 sky130_fd_sc_hd__and2_1 _07813_ (.A(_01437_),
    .B(_02353_),
    .X(_02354_));
 sky130_fd_sc_hd__buf_4 _07814_ (.A(_01405_),
    .X(_02355_));
 sky130_fd_sc_hd__a211o_1 _07815_ (.A1(_02346_),
    .A2(_02347_),
    .B1(_02354_),
    .C1(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__o211a_1 _07816_ (.A1(_01678_),
    .A2(_01973_),
    .B1(_01886_),
    .C1(_02356_),
    .X(_00265_));
 sky130_fd_sc_hd__xor2_4 _07817_ (.A(\_182_[23] ),
    .B(_01681_),
    .X(_02357_));
 sky130_fd_sc_hd__a21oi_2 _07818_ (.A1(_02350_),
    .A2(_02352_),
    .B1(_02349_),
    .Y(_02358_));
 sky130_fd_sc_hd__xnor2_4 _07819_ (.A(_02357_),
    .B(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__and2b_1 _07820_ (.A_N(_02336_),
    .B(_02337_),
    .X(_02360_));
 sky130_fd_sc_hd__xnor2_1 _07821_ (.A(_01657_),
    .B(_01608_),
    .Y(_02361_));
 sky130_fd_sc_hd__xnor2_2 _07822_ (.A(_01701_),
    .B(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__or2_1 _07823_ (.A(\_185_[23] ),
    .B(\_234_[23] ),
    .X(_02363_));
 sky130_fd_sc_hd__nand2_1 _07824_ (.A(\_185_[23] ),
    .B(\_234_[23] ),
    .Y(_02364_));
 sky130_fd_sc_hd__nand3_1 _07825_ (.A(_02362_),
    .B(_02363_),
    .C(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__a21o_1 _07826_ (.A1(_02363_),
    .A2(_02364_),
    .B1(_02362_),
    .X(_02366_));
 sky130_fd_sc_hd__nand2_1 _07827_ (.A(_02365_),
    .B(_02366_),
    .Y(_02367_));
 sky130_fd_sc_hd__a21oi_1 _07828_ (.A1(_02329_),
    .A2(_02331_),
    .B1(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__and3_1 _07829_ (.A(_02329_),
    .B(_02331_),
    .C(_02367_),
    .X(_02369_));
 sky130_fd_sc_hd__or2_1 _07830_ (.A(_02368_),
    .B(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__mux2_4 _07831_ (.A0(\_243_[23] ),
    .A1(\_240_[23] ),
    .S(_01681_),
    .X(_02371_));
 sky130_fd_sc_hd__xnor2_1 _07832_ (.A(_02370_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__nor3_1 _07833_ (.A(_02334_),
    .B(_02360_),
    .C(_02372_),
    .Y(_02373_));
 sky130_fd_sc_hd__o21ai_1 _07834_ (.A1(_02334_),
    .A2(_02360_),
    .B1(_02372_),
    .Y(_02374_));
 sky130_fd_sc_hd__and2b_1 _07835_ (.A_N(_02373_),
    .B(_02374_),
    .X(_02375_));
 sky130_fd_sc_hd__a21bo_1 _07836_ (.A1(_02341_),
    .A2(_02345_),
    .B1_N(_02339_),
    .X(_02376_));
 sky130_fd_sc_hd__nand2_1 _07837_ (.A(_02375_),
    .B(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__o211a_1 _07838_ (.A1(_02375_),
    .A2(_02376_),
    .B1(_02377_),
    .C1(_01523_),
    .X(_02378_));
 sky130_fd_sc_hd__a211o_1 _07839_ (.A1(_01856_),
    .A2(_02359_),
    .B1(_02378_),
    .C1(_02355_),
    .X(_02379_));
 sky130_fd_sc_hd__o211a_1 _07840_ (.A1(_01681_),
    .A2(_01973_),
    .B1(_01886_),
    .C1(_02379_),
    .X(_00266_));
 sky130_fd_sc_hd__buf_4 _07841_ (.A(_01437_),
    .X(_02380_));
 sky130_fd_sc_hd__and2b_1 _07842_ (.A_N(_02370_),
    .B(_02371_),
    .X(_02381_));
 sky130_fd_sc_hd__xnor2_2 _07843_ (.A(_01661_),
    .B(_01612_),
    .Y(_02382_));
 sky130_fd_sc_hd__xnor2_4 _07844_ (.A(_01704_),
    .B(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__or2_1 _07845_ (.A(\_185_[24] ),
    .B(\_234_[24] ),
    .X(_02384_));
 sky130_fd_sc_hd__nand2_1 _07846_ (.A(\_185_[24] ),
    .B(\_234_[24] ),
    .Y(_02385_));
 sky130_fd_sc_hd__nand3_1 _07847_ (.A(_02383_),
    .B(_02384_),
    .C(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__a21o_1 _07848_ (.A1(_02384_),
    .A2(_02385_),
    .B1(_02383_),
    .X(_02387_));
 sky130_fd_sc_hd__nand2_1 _07849_ (.A(_02386_),
    .B(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__a21oi_1 _07850_ (.A1(_02364_),
    .A2(_02365_),
    .B1(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__and3_1 _07851_ (.A(_02364_),
    .B(_02365_),
    .C(_02388_),
    .X(_02390_));
 sky130_fd_sc_hd__or2_1 _07852_ (.A(_02389_),
    .B(_02390_),
    .X(_02391_));
 sky130_fd_sc_hd__mux2_4 _07853_ (.A0(\_243_[24] ),
    .A1(\_240_[24] ),
    .S(_01684_),
    .X(_02392_));
 sky130_fd_sc_hd__xnor2_1 _07854_ (.A(_02391_),
    .B(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__o21ai_1 _07855_ (.A1(_02368_),
    .A2(_02381_),
    .B1(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__or3_1 _07856_ (.A(_02368_),
    .B(_02381_),
    .C(_02393_),
    .X(_02395_));
 sky130_fd_sc_hd__and2_1 _07857_ (.A(_02394_),
    .B(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__nand2_1 _07858_ (.A(_02341_),
    .B(_02375_),
    .Y(_02397_));
 sky130_fd_sc_hd__o221a_1 _07859_ (.A1(_02339_),
    .A2(_02373_),
    .B1(_02397_),
    .B2(_02344_),
    .C1(_02374_),
    .X(_02398_));
 sky130_fd_sc_hd__or2_1 _07860_ (.A(_02342_),
    .B(_02397_),
    .X(_02399_));
 sky130_fd_sc_hd__or2_1 _07861_ (.A(_02280_),
    .B(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__a211o_1 _07862_ (.A1(_02144_),
    .A2(_02147_),
    .B1(_02277_),
    .C1(_02399_),
    .X(_02401_));
 sky130_fd_sc_hd__and3_1 _07863_ (.A(_02398_),
    .B(_02400_),
    .C(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__xnor2_1 _07864_ (.A(_02396_),
    .B(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__clkbuf_4 _07865_ (.A(_01408_),
    .X(_02404_));
 sky130_fd_sc_hd__or2_1 _07866_ (.A(\_182_[24] ),
    .B(_01684_),
    .X(_02405_));
 sky130_fd_sc_hd__nand2_1 _07867_ (.A(\_182_[24] ),
    .B(_01684_),
    .Y(_02406_));
 sky130_fd_sc_hd__or4bb_1 _07868_ (.A(_02290_),
    .B(_02298_),
    .C_N(_02350_),
    .D_N(_02357_),
    .X(_02407_));
 sky130_fd_sc_hd__o21ba_1 _07869_ (.A1(\_182_[20] ),
    .A2(_01671_),
    .B1_N(_02285_),
    .X(_02408_));
 sky130_fd_sc_hd__o21a_1 _07870_ (.A1(_02351_),
    .A2(_02408_),
    .B1(_02297_),
    .X(_02409_));
 sky130_fd_sc_hd__or2_1 _07871_ (.A(\_182_[22] ),
    .B(_01678_),
    .X(_02410_));
 sky130_fd_sc_hd__o221a_1 _07872_ (.A1(\_182_[23] ),
    .A2(_01681_),
    .B1(_02349_),
    .B2(_02409_),
    .C1(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__a21oi_1 _07873_ (.A1(\_182_[23] ),
    .A2(_01681_),
    .B1(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__o31ai_2 _07874_ (.A1(_02172_),
    .A2(_02286_),
    .A3(_02407_),
    .B1(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__and3_1 _07875_ (.A(_02405_),
    .B(_02406_),
    .C(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__a21oi_1 _07876_ (.A1(_02405_),
    .A2(_02406_),
    .B1(_02413_),
    .Y(_02415_));
 sky130_fd_sc_hd__or2_2 _07877_ (.A(_02414_),
    .B(_02415_),
    .X(_02416_));
 sky130_fd_sc_hd__nand2_1 _07878_ (.A(_02404_),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__o211a_1 _07879_ (.A1(_02380_),
    .A2(_02403_),
    .B1(_02417_),
    .C1(_02202_),
    .X(_02418_));
 sky130_fd_sc_hd__a211o_1 _07880_ (.A1(_01684_),
    .A2(_01827_),
    .B1(_02178_),
    .C1(_02418_),
    .X(_00267_));
 sky130_fd_sc_hd__clkbuf_4 _07881_ (.A(_01480_),
    .X(_02419_));
 sky130_fd_sc_hd__and2b_1 _07882_ (.A_N(_02391_),
    .B(_02392_),
    .X(_02420_));
 sky130_fd_sc_hd__xnor2_2 _07883_ (.A(_01664_),
    .B(_01616_),
    .Y(_02421_));
 sky130_fd_sc_hd__xnor2_4 _07884_ (.A(_01707_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__or2_1 _07885_ (.A(\_185_[25] ),
    .B(\_234_[25] ),
    .X(_02423_));
 sky130_fd_sc_hd__nand2_1 _07886_ (.A(\_185_[25] ),
    .B(\_234_[25] ),
    .Y(_02424_));
 sky130_fd_sc_hd__nand3_1 _07887_ (.A(_02422_),
    .B(_02423_),
    .C(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__a21o_1 _07888_ (.A1(_02423_),
    .A2(_02424_),
    .B1(_02422_),
    .X(_02426_));
 sky130_fd_sc_hd__nand2_1 _07889_ (.A(_02425_),
    .B(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__a21oi_1 _07890_ (.A1(_02385_),
    .A2(_02386_),
    .B1(_02427_),
    .Y(_02428_));
 sky130_fd_sc_hd__and3_1 _07891_ (.A(_02385_),
    .B(_02386_),
    .C(_02427_),
    .X(_02429_));
 sky130_fd_sc_hd__or2_1 _07892_ (.A(_02428_),
    .B(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_4 _07893_ (.A0(\_243_[25] ),
    .A1(\_240_[25] ),
    .S(_01687_),
    .X(_02431_));
 sky130_fd_sc_hd__xnor2_1 _07894_ (.A(_02430_),
    .B(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__o21ai_1 _07895_ (.A1(_02389_),
    .A2(_02420_),
    .B1(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__inv_2 _07896_ (.A(_02433_),
    .Y(_02434_));
 sky130_fd_sc_hd__nor3_1 _07897_ (.A(_02389_),
    .B(_02420_),
    .C(_02432_),
    .Y(_02435_));
 sky130_fd_sc_hd__nor2_1 _07898_ (.A(_02434_),
    .B(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__inv_2 _07899_ (.A(_02396_),
    .Y(_02437_));
 sky130_fd_sc_hd__o21ai_1 _07900_ (.A1(_02437_),
    .A2(_02402_),
    .B1(_02394_),
    .Y(_02438_));
 sky130_fd_sc_hd__nand2_1 _07901_ (.A(_02436_),
    .B(_02438_),
    .Y(_02439_));
 sky130_fd_sc_hd__or2_1 _07902_ (.A(_02436_),
    .B(_02438_),
    .X(_02440_));
 sky130_fd_sc_hd__nand2_1 _07903_ (.A(\_182_[25] ),
    .B(_01687_),
    .Y(_02441_));
 sky130_fd_sc_hd__or2_1 _07904_ (.A(\_182_[25] ),
    .B(_01687_),
    .X(_02442_));
 sky130_fd_sc_hd__nand2_1 _07905_ (.A(_02441_),
    .B(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__a21oi_2 _07906_ (.A1(\_182_[24] ),
    .A2(_01684_),
    .B1(_02414_),
    .Y(_02444_));
 sky130_fd_sc_hd__xnor2_2 _07907_ (.A(_02443_),
    .B(_02444_),
    .Y(_02445_));
 sky130_fd_sc_hd__o21ai_2 _07908_ (.A1(_01778_),
    .A2(_02445_),
    .B1(_01412_),
    .Y(_02446_));
 sky130_fd_sc_hd__a31o_1 _07909_ (.A1(_01355_),
    .A2(_02439_),
    .A3(_02440_),
    .B1(_02446_),
    .X(_02447_));
 sky130_fd_sc_hd__o211a_1 _07910_ (.A1(_01687_),
    .A2(_01973_),
    .B1(_02419_),
    .C1(_02447_),
    .X(_00268_));
 sky130_fd_sc_hd__clkbuf_4 _07911_ (.A(_01421_),
    .X(_02448_));
 sky130_fd_sc_hd__and2b_1 _07912_ (.A_N(_02430_),
    .B(_02431_),
    .X(_02449_));
 sky130_fd_sc_hd__xnor2_2 _07913_ (.A(_01620_),
    .B(\_237_[0] ),
    .Y(_02450_));
 sky130_fd_sc_hd__xnor2_4 _07914_ (.A(_01667_),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__or2_1 _07915_ (.A(\_185_[26] ),
    .B(\_234_[26] ),
    .X(_02452_));
 sky130_fd_sc_hd__nand2_1 _07916_ (.A(\_185_[26] ),
    .B(\_234_[26] ),
    .Y(_02453_));
 sky130_fd_sc_hd__nand3_1 _07917_ (.A(_02451_),
    .B(_02452_),
    .C(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__a21o_1 _07918_ (.A1(_02452_),
    .A2(_02453_),
    .B1(_02451_),
    .X(_02455_));
 sky130_fd_sc_hd__nand2_1 _07919_ (.A(_02454_),
    .B(_02455_),
    .Y(_02456_));
 sky130_fd_sc_hd__a21oi_1 _07920_ (.A1(_02424_),
    .A2(_02425_),
    .B1(_02456_),
    .Y(_02457_));
 sky130_fd_sc_hd__and3_1 _07921_ (.A(_02424_),
    .B(_02425_),
    .C(_02456_),
    .X(_02458_));
 sky130_fd_sc_hd__or2_1 _07922_ (.A(_02457_),
    .B(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_4 _07923_ (.A0(\_243_[26] ),
    .A1(\_240_[26] ),
    .S(_01690_),
    .X(_02460_));
 sky130_fd_sc_hd__xnor2_1 _07924_ (.A(_02459_),
    .B(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__o21a_1 _07925_ (.A1(_02428_),
    .A2(_02449_),
    .B1(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__inv_2 _07926_ (.A(_02462_),
    .Y(_02463_));
 sky130_fd_sc_hd__or3_1 _07927_ (.A(_02428_),
    .B(_02449_),
    .C(_02461_),
    .X(_02464_));
 sky130_fd_sc_hd__and2_1 _07928_ (.A(_02463_),
    .B(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__nand2_1 _07929_ (.A(_02396_),
    .B(_02436_),
    .Y(_02466_));
 sky130_fd_sc_hd__nor2_1 _07930_ (.A(_02402_),
    .B(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__a21oi_1 _07931_ (.A1(_02394_),
    .A2(_02433_),
    .B1(_02435_),
    .Y(_02468_));
 sky130_fd_sc_hd__or3_1 _07932_ (.A(_02465_),
    .B(_02467_),
    .C(_02468_),
    .X(_02469_));
 sky130_fd_sc_hd__o21ai_1 _07933_ (.A1(_02467_),
    .A2(_02468_),
    .B1(_02465_),
    .Y(_02470_));
 sky130_fd_sc_hd__or2_1 _07934_ (.A(\_182_[26] ),
    .B(_01690_),
    .X(_02471_));
 sky130_fd_sc_hd__nand2_1 _07935_ (.A(\_182_[26] ),
    .B(_01690_),
    .Y(_02472_));
 sky130_fd_sc_hd__nand2_1 _07936_ (.A(_02471_),
    .B(_02472_),
    .Y(_02473_));
 sky130_fd_sc_hd__nor2_1 _07937_ (.A(\_182_[25] ),
    .B(_01687_),
    .Y(_02474_));
 sky130_fd_sc_hd__a21o_1 _07938_ (.A1(_02441_),
    .A2(_02444_),
    .B1(_02474_),
    .X(_02475_));
 sky130_fd_sc_hd__xnor2_2 _07939_ (.A(_02473_),
    .B(_02475_),
    .Y(_02476_));
 sky130_fd_sc_hd__o21ai_2 _07940_ (.A1(_01354_),
    .A2(_02476_),
    .B1(_01412_),
    .Y(_02477_));
 sky130_fd_sc_hd__a31o_1 _07941_ (.A1(_01355_),
    .A2(_02469_),
    .A3(_02470_),
    .B1(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__o211a_1 _07942_ (.A1(_01690_),
    .A2(_02448_),
    .B1(_02419_),
    .C1(_02478_),
    .X(_00269_));
 sky130_fd_sc_hd__nor2_1 _07943_ (.A(\_182_[27] ),
    .B(_01694_),
    .Y(_02479_));
 sky130_fd_sc_hd__nand2_1 _07944_ (.A(\_182_[27] ),
    .B(_01694_),
    .Y(_02480_));
 sky130_fd_sc_hd__or2b_1 _07945_ (.A(_02479_),
    .B_N(_02480_),
    .X(_02481_));
 sky130_fd_sc_hd__o21a_1 _07946_ (.A1(_02473_),
    .A2(_02475_),
    .B1(_02472_),
    .X(_02482_));
 sky130_fd_sc_hd__xor2_2 _07947_ (.A(_02481_),
    .B(_02482_),
    .X(_02483_));
 sky130_fd_sc_hd__and2b_1 _07948_ (.A_N(_02459_),
    .B(_02460_),
    .X(_02484_));
 sky130_fd_sc_hd__xnor2_2 _07949_ (.A(_01623_),
    .B(_01604_),
    .Y(_02485_));
 sky130_fd_sc_hd__xnor2_4 _07950_ (.A(_01671_),
    .B(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__or2_1 _07951_ (.A(\_185_[27] ),
    .B(\_234_[27] ),
    .X(_02487_));
 sky130_fd_sc_hd__nand2_1 _07952_ (.A(\_185_[27] ),
    .B(\_234_[27] ),
    .Y(_02488_));
 sky130_fd_sc_hd__nand3_1 _07953_ (.A(_02486_),
    .B(_02487_),
    .C(_02488_),
    .Y(_02489_));
 sky130_fd_sc_hd__a21o_1 _07954_ (.A1(_02487_),
    .A2(_02488_),
    .B1(_02486_),
    .X(_02490_));
 sky130_fd_sc_hd__nand2_1 _07955_ (.A(_02489_),
    .B(_02490_),
    .Y(_02491_));
 sky130_fd_sc_hd__a21oi_1 _07956_ (.A1(_02453_),
    .A2(_02454_),
    .B1(_02491_),
    .Y(_02492_));
 sky130_fd_sc_hd__and3_1 _07957_ (.A(_02453_),
    .B(_02454_),
    .C(_02491_),
    .X(_02493_));
 sky130_fd_sc_hd__or2_1 _07958_ (.A(_02492_),
    .B(_02493_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_4 _07959_ (.A0(\_243_[27] ),
    .A1(\_240_[27] ),
    .S(_01694_),
    .X(_02495_));
 sky130_fd_sc_hd__xnor2_1 _07960_ (.A(_02494_),
    .B(_02495_),
    .Y(_02496_));
 sky130_fd_sc_hd__nor3_1 _07961_ (.A(_02457_),
    .B(_02484_),
    .C(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__o21a_1 _07962_ (.A1(_02457_),
    .A2(_02484_),
    .B1(_02496_),
    .X(_02498_));
 sky130_fd_sc_hd__nor2_1 _07963_ (.A(_02497_),
    .B(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__and3_1 _07964_ (.A(_02463_),
    .B(_02470_),
    .C(_02499_),
    .X(_02500_));
 sky130_fd_sc_hd__a21oi_1 _07965_ (.A1(_02463_),
    .A2(_02470_),
    .B1(_02499_),
    .Y(_02501_));
 sky130_fd_sc_hd__o21a_1 _07966_ (.A1(_02500_),
    .A2(_02501_),
    .B1(_01354_),
    .X(_02502_));
 sky130_fd_sc_hd__a211o_1 _07967_ (.A1(_01856_),
    .A2(_02483_),
    .B1(_02502_),
    .C1(_02355_),
    .X(_02503_));
 sky130_fd_sc_hd__o211a_1 _07968_ (.A1(_01694_),
    .A2(_02448_),
    .B1(_02419_),
    .C1(_02503_),
    .X(_00270_));
 sky130_fd_sc_hd__and2b_1 _07969_ (.A_N(_02494_),
    .B(_02495_),
    .X(_02504_));
 sky130_fd_sc_hd__xnor2_2 _07970_ (.A(_01626_),
    .B(_01608_),
    .Y(_02505_));
 sky130_fd_sc_hd__xnor2_4 _07971_ (.A(_01675_),
    .B(_02505_),
    .Y(_02506_));
 sky130_fd_sc_hd__nand2_1 _07972_ (.A(\_185_[28] ),
    .B(\_234_[28] ),
    .Y(_02507_));
 sky130_fd_sc_hd__or2_1 _07973_ (.A(\_185_[28] ),
    .B(\_234_[28] ),
    .X(_02508_));
 sky130_fd_sc_hd__nand2_1 _07974_ (.A(_02507_),
    .B(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__xor2_1 _07975_ (.A(_02506_),
    .B(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__a21oi_1 _07976_ (.A1(_02488_),
    .A2(_02489_),
    .B1(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__and3_1 _07977_ (.A(_02488_),
    .B(_02489_),
    .C(_02510_),
    .X(_02512_));
 sky130_fd_sc_hd__or2_1 _07978_ (.A(_02511_),
    .B(_02512_),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_4 _07979_ (.A0(\_243_[28] ),
    .A1(\_240_[28] ),
    .S(_01698_),
    .X(_02514_));
 sky130_fd_sc_hd__xnor2_1 _07980_ (.A(_02513_),
    .B(_02514_),
    .Y(_02515_));
 sky130_fd_sc_hd__o21a_1 _07981_ (.A1(_02492_),
    .A2(_02504_),
    .B1(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__nor3_1 _07982_ (.A(_02492_),
    .B(_02504_),
    .C(_02515_),
    .Y(_02517_));
 sky130_fd_sc_hd__or2_1 _07983_ (.A(_02516_),
    .B(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__nand2_1 _07984_ (.A(_02465_),
    .B(_02499_),
    .Y(_02519_));
 sky130_fd_sc_hd__inv_2 _07985_ (.A(_02468_),
    .Y(_02520_));
 sky130_fd_sc_hd__inv_2 _07986_ (.A(_02498_),
    .Y(_02521_));
 sky130_fd_sc_hd__o221a_1 _07987_ (.A1(_02463_),
    .A2(_02497_),
    .B1(_02519_),
    .B2(_02520_),
    .C1(_02521_),
    .X(_02522_));
 sky130_fd_sc_hd__o31a_1 _07988_ (.A1(_02402_),
    .A2(_02466_),
    .A3(_02519_),
    .B1(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__and2_1 _07989_ (.A(_02518_),
    .B(_02523_),
    .X(_02524_));
 sky130_fd_sc_hd__nor2_1 _07990_ (.A(_02518_),
    .B(_02523_),
    .Y(_02525_));
 sky130_fd_sc_hd__nor2_1 _07991_ (.A(_02524_),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__or3_1 _07992_ (.A(_02474_),
    .B(_02473_),
    .C(_02481_),
    .X(_02527_));
 sky130_fd_sc_hd__and2b_1 _07993_ (.A_N(_02527_),
    .B(_02441_),
    .X(_02528_));
 sky130_fd_sc_hd__a21o_1 _07994_ (.A1(_02406_),
    .A2(_02441_),
    .B1(_02527_),
    .X(_02529_));
 sky130_fd_sc_hd__o211ai_1 _07995_ (.A1(_02472_),
    .A2(_02479_),
    .B1(_02480_),
    .C1(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__a21oi_2 _07996_ (.A1(_02414_),
    .A2(_02528_),
    .B1(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__nor2_1 _07997_ (.A(\_182_[28] ),
    .B(_01698_),
    .Y(_02532_));
 sky130_fd_sc_hd__nand2_1 _07998_ (.A(\_182_[28] ),
    .B(_01698_),
    .Y(_02533_));
 sky130_fd_sc_hd__or2b_1 _07999_ (.A(_02532_),
    .B_N(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__xnor2_2 _08000_ (.A(_02531_),
    .B(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__nand2_1 _08001_ (.A(_02404_),
    .B(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__o211a_1 _08002_ (.A1(_02380_),
    .A2(_02526_),
    .B1(_02536_),
    .C1(_02202_),
    .X(_02537_));
 sky130_fd_sc_hd__a211o_1 _08003_ (.A1(_01698_),
    .A2(_01827_),
    .B1(_02178_),
    .C1(_02537_),
    .X(_00271_));
 sky130_fd_sc_hd__and2b_1 _08004_ (.A_N(_02513_),
    .B(_02514_),
    .X(_02538_));
 sky130_fd_sc_hd__xnor2_2 _08005_ (.A(_01629_),
    .B(_01612_),
    .Y(_02539_));
 sky130_fd_sc_hd__xnor2_4 _08006_ (.A(_01678_),
    .B(_02539_),
    .Y(_02540_));
 sky130_fd_sc_hd__nand2_1 _08007_ (.A(\_185_[29] ),
    .B(\_234_[29] ),
    .Y(_02541_));
 sky130_fd_sc_hd__or2_1 _08008_ (.A(\_185_[29] ),
    .B(\_234_[29] ),
    .X(_02542_));
 sky130_fd_sc_hd__nand2_1 _08009_ (.A(_02541_),
    .B(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__xor2_1 _08010_ (.A(_02540_),
    .B(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__a21boi_1 _08011_ (.A1(_02506_),
    .A2(_02508_),
    .B1_N(_02507_),
    .Y(_02545_));
 sky130_fd_sc_hd__nor2_1 _08012_ (.A(_02544_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__and2_1 _08013_ (.A(_02544_),
    .B(_02545_),
    .X(_02547_));
 sky130_fd_sc_hd__or2_1 _08014_ (.A(_02546_),
    .B(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__mux2_4 _08015_ (.A0(\_243_[29] ),
    .A1(\_240_[29] ),
    .S(_01701_),
    .X(_02549_));
 sky130_fd_sc_hd__xnor2_1 _08016_ (.A(_02548_),
    .B(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__o21ai_1 _08017_ (.A1(_02511_),
    .A2(_02538_),
    .B1(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__inv_2 _08018_ (.A(_02551_),
    .Y(_02552_));
 sky130_fd_sc_hd__nor3_1 _08019_ (.A(_02511_),
    .B(_02538_),
    .C(_02550_),
    .Y(_02553_));
 sky130_fd_sc_hd__nor2_1 _08020_ (.A(_02552_),
    .B(_02553_),
    .Y(_02554_));
 sky130_fd_sc_hd__o21ai_1 _08021_ (.A1(_02516_),
    .A2(_02525_),
    .B1(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__o31a_1 _08022_ (.A1(_02516_),
    .A2(_02525_),
    .A3(_02554_),
    .B1(_01523_),
    .X(_02556_));
 sky130_fd_sc_hd__nor2_1 _08023_ (.A(\_182_[29] ),
    .B(_01701_),
    .Y(_02557_));
 sky130_fd_sc_hd__nand2_1 _08024_ (.A(\_182_[29] ),
    .B(_01701_),
    .Y(_02558_));
 sky130_fd_sc_hd__or2b_1 _08025_ (.A(_02557_),
    .B_N(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__o21a_1 _08026_ (.A1(_02531_),
    .A2(_02532_),
    .B1(_02533_),
    .X(_02560_));
 sky130_fd_sc_hd__xnor2_2 _08027_ (.A(_02559_),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__nor2_1 _08028_ (.A(_01778_),
    .B(_02561_),
    .Y(_02562_));
 sky130_fd_sc_hd__a211o_1 _08029_ (.A1(_02555_),
    .A2(_02556_),
    .B1(_02562_),
    .C1(_02355_),
    .X(_02563_));
 sky130_fd_sc_hd__o211a_1 _08030_ (.A1(_01701_),
    .A2(_02448_),
    .B1(_02419_),
    .C1(_02563_),
    .X(_00272_));
 sky130_fd_sc_hd__clkbuf_4 _08031_ (.A(_01406_),
    .X(_02564_));
 sky130_fd_sc_hd__nand2_1 _08032_ (.A(\_182_[30] ),
    .B(_01704_),
    .Y(_02565_));
 sky130_fd_sc_hd__or2_1 _08033_ (.A(\_182_[30] ),
    .B(_01704_),
    .X(_02566_));
 sky130_fd_sc_hd__nand2_1 _08034_ (.A(_02565_),
    .B(_02566_),
    .Y(_02567_));
 sky130_fd_sc_hd__o211a_1 _08035_ (.A1(_02531_),
    .A2(_02532_),
    .B1(_02533_),
    .C1(_02558_),
    .X(_02568_));
 sky130_fd_sc_hd__nor2_1 _08036_ (.A(_02557_),
    .B(_02568_),
    .Y(_02569_));
 sky130_fd_sc_hd__xnor2_2 _08037_ (.A(_02567_),
    .B(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__and2b_1 _08038_ (.A_N(_02548_),
    .B(_02549_),
    .X(_02571_));
 sky130_fd_sc_hd__xnor2_2 _08039_ (.A(_01632_),
    .B(_01616_),
    .Y(_02572_));
 sky130_fd_sc_hd__xnor2_4 _08040_ (.A(_01681_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__nor2_1 _08041_ (.A(\_185_[30] ),
    .B(\_234_[30] ),
    .Y(_02574_));
 sky130_fd_sc_hd__and2_1 _08042_ (.A(\_185_[30] ),
    .B(\_234_[30] ),
    .X(_02575_));
 sky130_fd_sc_hd__nor2_1 _08043_ (.A(_02574_),
    .B(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__xnor2_1 _08044_ (.A(_02573_),
    .B(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__a21bo_1 _08045_ (.A1(_02540_),
    .A2(_02542_),
    .B1_N(_02541_),
    .X(_02578_));
 sky130_fd_sc_hd__and2b_1 _08046_ (.A_N(_02577_),
    .B(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__or2b_1 _08047_ (.A(_02578_),
    .B_N(_02577_),
    .X(_02580_));
 sky130_fd_sc_hd__or2b_1 _08048_ (.A(_02579_),
    .B_N(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_4 _08049_ (.A0(\_243_[30] ),
    .A1(\_240_[30] ),
    .S(_01704_),
    .X(_02582_));
 sky130_fd_sc_hd__xnor2_1 _08050_ (.A(_02581_),
    .B(_02582_),
    .Y(_02583_));
 sky130_fd_sc_hd__o21a_1 _08051_ (.A1(_02546_),
    .A2(_02571_),
    .B1(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__nor3_1 _08052_ (.A(_02546_),
    .B(_02571_),
    .C(_02583_),
    .Y(_02585_));
 sky130_fd_sc_hd__nor2_1 _08053_ (.A(_02584_),
    .B(_02585_),
    .Y(_02586_));
 sky130_fd_sc_hd__o21bai_1 _08054_ (.A1(_02516_),
    .A2(_02552_),
    .B1_N(_02553_),
    .Y(_02587_));
 sky130_fd_sc_hd__o41a_1 _08055_ (.A1(_02518_),
    .A2(_02523_),
    .A3(_02552_),
    .A4(_02553_),
    .B1(_02587_),
    .X(_02588_));
 sky130_fd_sc_hd__xnor2_1 _08056_ (.A(_02586_),
    .B(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__or2_1 _08057_ (.A(_01408_),
    .B(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__o211a_1 _08058_ (.A1(_01520_),
    .A2(_02570_),
    .B1(_02590_),
    .C1(_02202_),
    .X(_02591_));
 sky130_fd_sc_hd__a211o_1 _08059_ (.A1(_01704_),
    .A2(_02564_),
    .B1(_02178_),
    .C1(_02591_),
    .X(_00273_));
 sky130_fd_sc_hd__o21bai_1 _08060_ (.A1(_02585_),
    .A2(_02588_),
    .B1_N(_02584_),
    .Y(_02592_));
 sky130_fd_sc_hd__a21oi_1 _08061_ (.A1(_02580_),
    .A2(_02582_),
    .B1(_02579_),
    .Y(_02593_));
 sky130_fd_sc_hd__xnor2_1 _08062_ (.A(_01635_),
    .B(_01620_),
    .Y(_02594_));
 sky130_fd_sc_hd__xnor2_2 _08063_ (.A(_01684_),
    .B(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__mux2_2 _08064_ (.A0(\_243_[31] ),
    .A1(\_240_[31] ),
    .S(_01707_),
    .X(_02596_));
 sky130_fd_sc_hd__xor2_4 _08065_ (.A(\_185_[31] ),
    .B(_02596_),
    .X(_02597_));
 sky130_fd_sc_hd__xnor2_4 _08066_ (.A(_02595_),
    .B(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__a21o_1 _08067_ (.A1(_02573_),
    .A2(_02576_),
    .B1(_02575_),
    .X(_02599_));
 sky130_fd_sc_hd__xnor2_1 _08068_ (.A(\_234_[31] ),
    .B(_02599_),
    .Y(_02600_));
 sky130_fd_sc_hd__xnor2_1 _08069_ (.A(_02598_),
    .B(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__xnor2_1 _08070_ (.A(_02593_),
    .B(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__xnor2_1 _08071_ (.A(_02592_),
    .B(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hd__o31a_1 _08072_ (.A1(_02557_),
    .A2(_02567_),
    .A3(_02568_),
    .B1(_02565_),
    .X(_02604_));
 sky130_fd_sc_hd__xnor2_1 _08073_ (.A(\_182_[31] ),
    .B(_01707_),
    .Y(_02605_));
 sky130_fd_sc_hd__xnor2_2 _08074_ (.A(_02604_),
    .B(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__nor2_1 _08075_ (.A(_01778_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__a211o_1 _08076_ (.A1(_01355_),
    .A2(_02603_),
    .B1(_02607_),
    .C1(_02355_),
    .X(_02608_));
 sky130_fd_sc_hd__o211a_1 _08077_ (.A1(_01707_),
    .A2(_02448_),
    .B1(_02419_),
    .C1(_02608_),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _08078_ (.A0(\_167_[0] ),
    .A1(\_231_[0] ),
    .S(_01672_),
    .X(_02609_));
 sky130_fd_sc_hd__or2_1 _08079_ (.A(_01670_),
    .B(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__o211a_1 _08080_ (.A1(\_234_[0] ),
    .A2(_02448_),
    .B1(_02419_),
    .C1(_02610_),
    .X(_00275_));
 sky130_fd_sc_hd__clkbuf_4 _08081_ (.A(_01437_),
    .X(_02611_));
 sky130_fd_sc_hd__or2_1 _08082_ (.A(\_167_[1] ),
    .B(_01646_),
    .X(_02612_));
 sky130_fd_sc_hd__o211a_1 _08083_ (.A1(\_231_[1] ),
    .A2(_02611_),
    .B1(_01695_),
    .C1(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__a211o_1 _08084_ (.A1(\_234_[1] ),
    .A2(_02564_),
    .B1(_02178_),
    .C1(_02613_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _08085_ (.A0(\_167_[2] ),
    .A1(\_231_[2] ),
    .S(_01672_),
    .X(_02614_));
 sky130_fd_sc_hd__or2_1 _08086_ (.A(_01670_),
    .B(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__o211a_1 _08087_ (.A1(\_234_[2] ),
    .A2(_02448_),
    .B1(_02419_),
    .C1(_02615_),
    .X(_00277_));
 sky130_fd_sc_hd__clkbuf_2 _08088_ (.A(_01339_),
    .X(_02616_));
 sky130_fd_sc_hd__or2_1 _08089_ (.A(\_167_[3] ),
    .B(_02616_),
    .X(_02617_));
 sky130_fd_sc_hd__o211a_1 _08090_ (.A1(\_231_[3] ),
    .A2(_02611_),
    .B1(_01695_),
    .C1(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__a211o_1 _08091_ (.A1(\_234_[3] ),
    .A2(_02564_),
    .B1(_02178_),
    .C1(_02618_),
    .X(_00278_));
 sky130_fd_sc_hd__or2_1 _08092_ (.A(\_167_[4] ),
    .B(_02616_),
    .X(_02619_));
 sky130_fd_sc_hd__o211a_1 _08093_ (.A1(\_231_[4] ),
    .A2(_02611_),
    .B1(_01695_),
    .C1(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__a211o_1 _08094_ (.A1(\_234_[4] ),
    .A2(_02564_),
    .B1(_02178_),
    .C1(_02620_),
    .X(_00279_));
 sky130_fd_sc_hd__or2_1 _08095_ (.A(\_167_[5] ),
    .B(_02616_),
    .X(_02621_));
 sky130_fd_sc_hd__o211a_1 _08096_ (.A1(\_231_[5] ),
    .A2(_02611_),
    .B1(_01695_),
    .C1(_02621_),
    .X(_02622_));
 sky130_fd_sc_hd__a211o_1 _08097_ (.A1(\_234_[5] ),
    .A2(_02564_),
    .B1(_02178_),
    .C1(_02622_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _08098_ (.A0(\_167_[6] ),
    .A1(\_231_[6] ),
    .S(_01672_),
    .X(_02623_));
 sky130_fd_sc_hd__or2_1 _08099_ (.A(_01670_),
    .B(_02623_),
    .X(_02624_));
 sky130_fd_sc_hd__o211a_1 _08100_ (.A1(\_234_[6] ),
    .A2(_02448_),
    .B1(_02419_),
    .C1(_02624_),
    .X(_00281_));
 sky130_fd_sc_hd__clkbuf_2 _08101_ (.A(_01405_),
    .X(_02625_));
 sky130_fd_sc_hd__buf_4 _08102_ (.A(_01518_),
    .X(_02626_));
 sky130_fd_sc_hd__mux2_1 _08103_ (.A0(\_167_[7] ),
    .A1(\_231_[7] ),
    .S(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__or2_1 _08104_ (.A(_02625_),
    .B(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__o211a_1 _08105_ (.A1(\_234_[7] ),
    .A2(_02448_),
    .B1(_02419_),
    .C1(_02628_),
    .X(_00282_));
 sky130_fd_sc_hd__clkbuf_4 _08106_ (.A(_01435_),
    .X(_02629_));
 sky130_fd_sc_hd__or2_1 _08107_ (.A(\_167_[8] ),
    .B(_02616_),
    .X(_02630_));
 sky130_fd_sc_hd__o211a_1 _08108_ (.A1(\_231_[8] ),
    .A2(_02611_),
    .B1(_01695_),
    .C1(_02630_),
    .X(_02631_));
 sky130_fd_sc_hd__a211o_1 _08109_ (.A1(\_234_[8] ),
    .A2(_02564_),
    .B1(_02629_),
    .C1(_02631_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _08110_ (.A0(\_167_[9] ),
    .A1(\_231_[9] ),
    .S(_02626_),
    .X(_02632_));
 sky130_fd_sc_hd__or2_1 _08111_ (.A(_02625_),
    .B(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__o211a_1 _08112_ (.A1(\_234_[9] ),
    .A2(_02448_),
    .B1(_02419_),
    .C1(_02633_),
    .X(_00284_));
 sky130_fd_sc_hd__or2_1 _08113_ (.A(\_167_[10] ),
    .B(_02616_),
    .X(_02634_));
 sky130_fd_sc_hd__o211a_1 _08114_ (.A1(\_231_[10] ),
    .A2(_02611_),
    .B1(_01695_),
    .C1(_02634_),
    .X(_02635_));
 sky130_fd_sc_hd__a211o_1 _08115_ (.A1(\_234_[10] ),
    .A2(_02564_),
    .B1(_02629_),
    .C1(_02635_),
    .X(_00285_));
 sky130_fd_sc_hd__clkbuf_4 _08116_ (.A(_01480_),
    .X(_02636_));
 sky130_fd_sc_hd__mux2_1 _08117_ (.A0(\_167_[11] ),
    .A1(\_231_[11] ),
    .S(_02626_),
    .X(_02637_));
 sky130_fd_sc_hd__or2_1 _08118_ (.A(_02625_),
    .B(_02637_),
    .X(_02638_));
 sky130_fd_sc_hd__o211a_1 _08119_ (.A1(\_234_[11] ),
    .A2(_02448_),
    .B1(_02636_),
    .C1(_02638_),
    .X(_00286_));
 sky130_fd_sc_hd__or2_1 _08120_ (.A(\_167_[12] ),
    .B(_02616_),
    .X(_02639_));
 sky130_fd_sc_hd__o211a_1 _08121_ (.A1(\_231_[12] ),
    .A2(_02611_),
    .B1(_01695_),
    .C1(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__a211o_1 _08122_ (.A1(\_234_[12] ),
    .A2(_02564_),
    .B1(_02629_),
    .C1(_02640_),
    .X(_00287_));
 sky130_fd_sc_hd__clkbuf_4 _08123_ (.A(_01420_),
    .X(_02641_));
 sky130_fd_sc_hd__or2_1 _08124_ (.A(\_167_[13] ),
    .B(_02616_),
    .X(_02642_));
 sky130_fd_sc_hd__o211a_1 _08125_ (.A1(\_231_[13] ),
    .A2(_02611_),
    .B1(_02641_),
    .C1(_02642_),
    .X(_02643_));
 sky130_fd_sc_hd__a211o_1 _08126_ (.A1(\_234_[13] ),
    .A2(_02564_),
    .B1(_02629_),
    .C1(_02643_),
    .X(_00288_));
 sky130_fd_sc_hd__or2_1 _08127_ (.A(\_167_[14] ),
    .B(_02616_),
    .X(_02644_));
 sky130_fd_sc_hd__o211a_1 _08128_ (.A1(\_231_[14] ),
    .A2(_02611_),
    .B1(_02641_),
    .C1(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__a211o_1 _08129_ (.A1(\_234_[14] ),
    .A2(_02564_),
    .B1(_02629_),
    .C1(_02645_),
    .X(_00289_));
 sky130_fd_sc_hd__clkbuf_4 _08130_ (.A(_01406_),
    .X(_02646_));
 sky130_fd_sc_hd__or2_1 _08131_ (.A(\_167_[15] ),
    .B(_02616_),
    .X(_02647_));
 sky130_fd_sc_hd__o211a_1 _08132_ (.A1(\_231_[15] ),
    .A2(_02611_),
    .B1(_02641_),
    .C1(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__a211o_1 _08133_ (.A1(\_234_[15] ),
    .A2(_02646_),
    .B1(_02629_),
    .C1(_02648_),
    .X(_00290_));
 sky130_fd_sc_hd__clkbuf_4 _08134_ (.A(_01437_),
    .X(_02649_));
 sky130_fd_sc_hd__or2_1 _08135_ (.A(\_167_[16] ),
    .B(_02616_),
    .X(_02650_));
 sky130_fd_sc_hd__o211a_1 _08136_ (.A1(\_231_[16] ),
    .A2(_02649_),
    .B1(_02641_),
    .C1(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__a211o_1 _08137_ (.A1(\_234_[16] ),
    .A2(_02646_),
    .B1(_02629_),
    .C1(_02651_),
    .X(_00291_));
 sky130_fd_sc_hd__clkbuf_2 _08138_ (.A(_01339_),
    .X(_02652_));
 sky130_fd_sc_hd__or2_1 _08139_ (.A(\_167_[17] ),
    .B(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__o211a_1 _08140_ (.A1(\_231_[17] ),
    .A2(_02649_),
    .B1(_02641_),
    .C1(_02653_),
    .X(_02654_));
 sky130_fd_sc_hd__a211o_1 _08141_ (.A1(\_234_[17] ),
    .A2(_02646_),
    .B1(_02629_),
    .C1(_02654_),
    .X(_00292_));
 sky130_fd_sc_hd__or2_1 _08142_ (.A(\_167_[18] ),
    .B(_02652_),
    .X(_02655_));
 sky130_fd_sc_hd__o211a_1 _08143_ (.A1(\_231_[18] ),
    .A2(_02649_),
    .B1(_02641_),
    .C1(_02655_),
    .X(_02656_));
 sky130_fd_sc_hd__a211o_1 _08144_ (.A1(\_234_[18] ),
    .A2(_02646_),
    .B1(_02629_),
    .C1(_02656_),
    .X(_00293_));
 sky130_fd_sc_hd__or2_1 _08145_ (.A(\_167_[19] ),
    .B(_02652_),
    .X(_02657_));
 sky130_fd_sc_hd__o211a_1 _08146_ (.A1(\_231_[19] ),
    .A2(_02649_),
    .B1(_02641_),
    .C1(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__a211o_1 _08147_ (.A1(\_234_[19] ),
    .A2(_02646_),
    .B1(_02629_),
    .C1(_02658_),
    .X(_00294_));
 sky130_fd_sc_hd__clkbuf_4 _08148_ (.A(_01421_),
    .X(_02659_));
 sky130_fd_sc_hd__mux2_1 _08149_ (.A0(\_167_[20] ),
    .A1(\_231_[20] ),
    .S(_02626_),
    .X(_02660_));
 sky130_fd_sc_hd__or2_1 _08150_ (.A(_02625_),
    .B(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__o211a_1 _08151_ (.A1(\_234_[20] ),
    .A2(_02659_),
    .B1(_02636_),
    .C1(_02661_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _08152_ (.A0(\_167_[21] ),
    .A1(\_231_[21] ),
    .S(_02626_),
    .X(_02662_));
 sky130_fd_sc_hd__or2_1 _08153_ (.A(_02625_),
    .B(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__o211a_1 _08154_ (.A1(\_234_[21] ),
    .A2(_02659_),
    .B1(_02636_),
    .C1(_02663_),
    .X(_00296_));
 sky130_fd_sc_hd__clkbuf_4 _08155_ (.A(_01435_),
    .X(_02664_));
 sky130_fd_sc_hd__or2_1 _08156_ (.A(\_167_[22] ),
    .B(_02652_),
    .X(_02665_));
 sky130_fd_sc_hd__o211a_1 _08157_ (.A1(\_231_[22] ),
    .A2(_02649_),
    .B1(_02641_),
    .C1(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__a211o_1 _08158_ (.A1(\_234_[22] ),
    .A2(_02646_),
    .B1(_02664_),
    .C1(_02666_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _08159_ (.A0(\_167_[23] ),
    .A1(\_231_[23] ),
    .S(_02626_),
    .X(_02667_));
 sky130_fd_sc_hd__or2_1 _08160_ (.A(_02625_),
    .B(_02667_),
    .X(_02668_));
 sky130_fd_sc_hd__o211a_1 _08161_ (.A1(\_234_[23] ),
    .A2(_02659_),
    .B1(_02636_),
    .C1(_02668_),
    .X(_00298_));
 sky130_fd_sc_hd__or2_1 _08162_ (.A(\_167_[24] ),
    .B(_02652_),
    .X(_02669_));
 sky130_fd_sc_hd__o211a_1 _08163_ (.A1(\_231_[24] ),
    .A2(_02649_),
    .B1(_02641_),
    .C1(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__a211o_1 _08164_ (.A1(\_234_[24] ),
    .A2(_02646_),
    .B1(_02664_),
    .C1(_02670_),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _08165_ (.A0(\_167_[25] ),
    .A1(\_231_[25] ),
    .S(_02626_),
    .X(_02671_));
 sky130_fd_sc_hd__or2_1 _08166_ (.A(_02625_),
    .B(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__o211a_1 _08167_ (.A1(\_234_[25] ),
    .A2(_02659_),
    .B1(_02636_),
    .C1(_02672_),
    .X(_00300_));
 sky130_fd_sc_hd__or2_1 _08168_ (.A(\_167_[26] ),
    .B(_02652_),
    .X(_02673_));
 sky130_fd_sc_hd__o211a_1 _08169_ (.A1(\_231_[26] ),
    .A2(_02649_),
    .B1(_02641_),
    .C1(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__a211o_1 _08170_ (.A1(\_234_[26] ),
    .A2(_02646_),
    .B1(_02664_),
    .C1(_02674_),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _08171_ (.A0(\_167_[27] ),
    .A1(\_231_[27] ),
    .S(_02626_),
    .X(_02675_));
 sky130_fd_sc_hd__or2_1 _08172_ (.A(_02625_),
    .B(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__o211a_1 _08173_ (.A1(\_234_[27] ),
    .A2(_02659_),
    .B1(_02636_),
    .C1(_02676_),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _08174_ (.A0(\_167_[28] ),
    .A1(\_231_[28] ),
    .S(_02626_),
    .X(_02677_));
 sky130_fd_sc_hd__or2_1 _08175_ (.A(_02625_),
    .B(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__o211a_1 _08176_ (.A1(\_234_[28] ),
    .A2(_02659_),
    .B1(_02636_),
    .C1(_02678_),
    .X(_00303_));
 sky130_fd_sc_hd__clkbuf_4 _08177_ (.A(_01420_),
    .X(_02679_));
 sky130_fd_sc_hd__or2_1 _08178_ (.A(\_167_[29] ),
    .B(_02652_),
    .X(_02680_));
 sky130_fd_sc_hd__o211a_1 _08179_ (.A1(\_231_[29] ),
    .A2(_02649_),
    .B1(_02679_),
    .C1(_02680_),
    .X(_02681_));
 sky130_fd_sc_hd__a211o_1 _08180_ (.A1(\_234_[29] ),
    .A2(_02646_),
    .B1(_02664_),
    .C1(_02681_),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _08181_ (.A0(\_167_[30] ),
    .A1(\_231_[30] ),
    .S(_02626_),
    .X(_02682_));
 sky130_fd_sc_hd__or2_1 _08182_ (.A(_02625_),
    .B(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__o211a_1 _08183_ (.A1(\_234_[30] ),
    .A2(_02659_),
    .B1(_02636_),
    .C1(_02683_),
    .X(_00305_));
 sky130_fd_sc_hd__or2_1 _08184_ (.A(\_167_[31] ),
    .B(_02652_),
    .X(_02684_));
 sky130_fd_sc_hd__o211a_1 _08185_ (.A1(\_231_[31] ),
    .A2(_02649_),
    .B1(_02679_),
    .C1(_02684_),
    .X(_02685_));
 sky130_fd_sc_hd__a211o_1 _08186_ (.A1(\_234_[31] ),
    .A2(_02646_),
    .B1(_02664_),
    .C1(_02685_),
    .X(_00306_));
 sky130_fd_sc_hd__buf_2 _08187_ (.A(_01405_),
    .X(_02686_));
 sky130_fd_sc_hd__buf_4 _08188_ (.A(_01518_),
    .X(_02687_));
 sky130_fd_sc_hd__mux2_1 _08189_ (.A0(\_164_[0] ),
    .A1(\_228_[0] ),
    .S(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__or2_1 _08190_ (.A(_02686_),
    .B(_02688_),
    .X(_02689_));
 sky130_fd_sc_hd__o211a_1 _08191_ (.A1(\_231_[0] ),
    .A2(_02659_),
    .B1(_02636_),
    .C1(_02689_),
    .X(_00307_));
 sky130_fd_sc_hd__clkbuf_4 _08192_ (.A(_01406_),
    .X(_02690_));
 sky130_fd_sc_hd__or2_1 _08193_ (.A(\_164_[1] ),
    .B(_02652_),
    .X(_02691_));
 sky130_fd_sc_hd__o211a_1 _08194_ (.A1(\_228_[1] ),
    .A2(_02649_),
    .B1(_02679_),
    .C1(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__a211o_1 _08195_ (.A1(\_231_[1] ),
    .A2(_02690_),
    .B1(_02664_),
    .C1(_02692_),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _08196_ (.A0(\_164_[2] ),
    .A1(\_228_[2] ),
    .S(_02687_),
    .X(_02693_));
 sky130_fd_sc_hd__or2_1 _08197_ (.A(_02686_),
    .B(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__o211a_1 _08198_ (.A1(\_231_[2] ),
    .A2(_02659_),
    .B1(_02636_),
    .C1(_02694_),
    .X(_00309_));
 sky130_fd_sc_hd__clkbuf_4 _08199_ (.A(_01480_),
    .X(_02695_));
 sky130_fd_sc_hd__mux2_1 _08200_ (.A0(\_164_[3] ),
    .A1(\_228_[3] ),
    .S(_02687_),
    .X(_02696_));
 sky130_fd_sc_hd__or2_1 _08201_ (.A(_02686_),
    .B(_02696_),
    .X(_02697_));
 sky130_fd_sc_hd__o211a_1 _08202_ (.A1(\_231_[3] ),
    .A2(_02659_),
    .B1(_02695_),
    .C1(_02697_),
    .X(_00310_));
 sky130_fd_sc_hd__clkbuf_4 _08203_ (.A(_01437_),
    .X(_02698_));
 sky130_fd_sc_hd__or2_1 _08204_ (.A(\_164_[4] ),
    .B(_02652_),
    .X(_02699_));
 sky130_fd_sc_hd__o211a_1 _08205_ (.A1(\_228_[4] ),
    .A2(_02698_),
    .B1(_02679_),
    .C1(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__a211o_1 _08206_ (.A1(\_231_[4] ),
    .A2(_02690_),
    .B1(_02664_),
    .C1(_02700_),
    .X(_00311_));
 sky130_fd_sc_hd__clkbuf_2 _08207_ (.A(_01339_),
    .X(_02701_));
 sky130_fd_sc_hd__or2_1 _08208_ (.A(\_164_[5] ),
    .B(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__o211a_1 _08209_ (.A1(\_228_[5] ),
    .A2(_02698_),
    .B1(_02679_),
    .C1(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__a211o_1 _08210_ (.A1(\_231_[5] ),
    .A2(_02690_),
    .B1(_02664_),
    .C1(_02703_),
    .X(_00312_));
 sky130_fd_sc_hd__or2_1 _08211_ (.A(\_164_[6] ),
    .B(_02701_),
    .X(_02704_));
 sky130_fd_sc_hd__o211a_1 _08212_ (.A1(\_228_[6] ),
    .A2(_02698_),
    .B1(_02679_),
    .C1(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__a211o_1 _08213_ (.A1(\_231_[6] ),
    .A2(_02690_),
    .B1(_02664_),
    .C1(_02705_),
    .X(_00313_));
 sky130_fd_sc_hd__buf_2 _08214_ (.A(_01799_),
    .X(_02706_));
 sky130_fd_sc_hd__mux2_1 _08215_ (.A0(\_164_[7] ),
    .A1(\_228_[7] ),
    .S(_02687_),
    .X(_02707_));
 sky130_fd_sc_hd__or2_1 _08216_ (.A(_02686_),
    .B(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__o211a_1 _08217_ (.A1(\_231_[7] ),
    .A2(_02706_),
    .B1(_02695_),
    .C1(_02708_),
    .X(_00314_));
 sky130_fd_sc_hd__or2_1 _08218_ (.A(\_164_[8] ),
    .B(_02701_),
    .X(_02709_));
 sky130_fd_sc_hd__o211a_1 _08219_ (.A1(\_228_[8] ),
    .A2(_02698_),
    .B1(_02679_),
    .C1(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__a211o_1 _08220_ (.A1(\_231_[8] ),
    .A2(_02690_),
    .B1(_02664_),
    .C1(_02710_),
    .X(_00315_));
 sky130_fd_sc_hd__buf_4 _08221_ (.A(_01417_),
    .X(_02711_));
 sky130_fd_sc_hd__clkbuf_4 _08222_ (.A(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__or2_1 _08223_ (.A(\_164_[9] ),
    .B(_02701_),
    .X(_02713_));
 sky130_fd_sc_hd__o211a_1 _08224_ (.A1(\_228_[9] ),
    .A2(_02698_),
    .B1(_02679_),
    .C1(_02713_),
    .X(_02714_));
 sky130_fd_sc_hd__a211o_1 _08225_ (.A1(\_231_[9] ),
    .A2(_02690_),
    .B1(_02712_),
    .C1(_02714_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _08226_ (.A0(\_164_[10] ),
    .A1(\_228_[10] ),
    .S(_02687_),
    .X(_02715_));
 sky130_fd_sc_hd__or2_1 _08227_ (.A(_02686_),
    .B(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__o211a_1 _08228_ (.A1(\_231_[10] ),
    .A2(_02706_),
    .B1(_02695_),
    .C1(_02716_),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _08229_ (.A0(\_164_[11] ),
    .A1(\_228_[11] ),
    .S(_02687_),
    .X(_02717_));
 sky130_fd_sc_hd__or2_1 _08230_ (.A(_02686_),
    .B(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__o211a_1 _08231_ (.A1(\_231_[11] ),
    .A2(_02706_),
    .B1(_02695_),
    .C1(_02718_),
    .X(_00318_));
 sky130_fd_sc_hd__or2_1 _08232_ (.A(\_164_[12] ),
    .B(_02701_),
    .X(_02719_));
 sky130_fd_sc_hd__o211a_1 _08233_ (.A1(\_228_[12] ),
    .A2(_02698_),
    .B1(_02679_),
    .C1(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__a211o_1 _08234_ (.A1(\_231_[12] ),
    .A2(_02690_),
    .B1(_02712_),
    .C1(_02720_),
    .X(_00319_));
 sky130_fd_sc_hd__or2_1 _08235_ (.A(\_164_[13] ),
    .B(_02701_),
    .X(_02721_));
 sky130_fd_sc_hd__o211a_1 _08236_ (.A1(\_228_[13] ),
    .A2(_02698_),
    .B1(_02679_),
    .C1(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__a211o_1 _08237_ (.A1(\_231_[13] ),
    .A2(_02690_),
    .B1(_02712_),
    .C1(_02722_),
    .X(_00320_));
 sky130_fd_sc_hd__clkbuf_4 _08238_ (.A(_01420_),
    .X(_02723_));
 sky130_fd_sc_hd__or2_1 _08239_ (.A(\_164_[14] ),
    .B(_02701_),
    .X(_02724_));
 sky130_fd_sc_hd__o211a_1 _08240_ (.A1(\_228_[14] ),
    .A2(_02698_),
    .B1(_02723_),
    .C1(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__a211o_1 _08241_ (.A1(\_231_[14] ),
    .A2(_02690_),
    .B1(_02712_),
    .C1(_02725_),
    .X(_00321_));
 sky130_fd_sc_hd__or2_1 _08242_ (.A(\_164_[15] ),
    .B(_02701_),
    .X(_02726_));
 sky130_fd_sc_hd__o211a_1 _08243_ (.A1(\_228_[15] ),
    .A2(_02698_),
    .B1(_02723_),
    .C1(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__a211o_1 _08244_ (.A1(\_231_[15] ),
    .A2(_02690_),
    .B1(_02712_),
    .C1(_02727_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _08245_ (.A0(\_164_[16] ),
    .A1(\_228_[16] ),
    .S(_02687_),
    .X(_02728_));
 sky130_fd_sc_hd__or2_1 _08246_ (.A(_02686_),
    .B(_02728_),
    .X(_02729_));
 sky130_fd_sc_hd__o211a_1 _08247_ (.A1(\_231_[16] ),
    .A2(_02706_),
    .B1(_02695_),
    .C1(_02729_),
    .X(_00323_));
 sky130_fd_sc_hd__clkbuf_4 _08248_ (.A(_01406_),
    .X(_02730_));
 sky130_fd_sc_hd__or2_1 _08249_ (.A(\_164_[17] ),
    .B(_02701_),
    .X(_02731_));
 sky130_fd_sc_hd__o211a_1 _08250_ (.A1(\_228_[17] ),
    .A2(_02698_),
    .B1(_02723_),
    .C1(_02731_),
    .X(_02732_));
 sky130_fd_sc_hd__a211o_1 _08251_ (.A1(\_231_[17] ),
    .A2(_02730_),
    .B1(_02712_),
    .C1(_02732_),
    .X(_00324_));
 sky130_fd_sc_hd__clkbuf_4 _08252_ (.A(_01437_),
    .X(_02733_));
 sky130_fd_sc_hd__or2_1 _08253_ (.A(\_164_[18] ),
    .B(_02701_),
    .X(_02734_));
 sky130_fd_sc_hd__o211a_1 _08254_ (.A1(\_228_[18] ),
    .A2(_02733_),
    .B1(_02723_),
    .C1(_02734_),
    .X(_02735_));
 sky130_fd_sc_hd__a211o_1 _08255_ (.A1(\_231_[18] ),
    .A2(_02730_),
    .B1(_02712_),
    .C1(_02735_),
    .X(_00325_));
 sky130_fd_sc_hd__buf_2 _08256_ (.A(_01339_),
    .X(_02736_));
 sky130_fd_sc_hd__or2_1 _08257_ (.A(\_164_[19] ),
    .B(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__o211a_1 _08258_ (.A1(\_228_[19] ),
    .A2(_02733_),
    .B1(_02723_),
    .C1(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__a211o_1 _08259_ (.A1(\_231_[19] ),
    .A2(_02730_),
    .B1(_02712_),
    .C1(_02738_),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _08260_ (.A0(\_164_[20] ),
    .A1(\_228_[20] ),
    .S(_02687_),
    .X(_02739_));
 sky130_fd_sc_hd__or2_1 _08261_ (.A(_02686_),
    .B(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__o211a_1 _08262_ (.A1(\_231_[20] ),
    .A2(_02706_),
    .B1(_02695_),
    .C1(_02740_),
    .X(_00327_));
 sky130_fd_sc_hd__or2_1 _08263_ (.A(\_164_[21] ),
    .B(_02736_),
    .X(_02741_));
 sky130_fd_sc_hd__o211a_1 _08264_ (.A1(\_228_[21] ),
    .A2(_02733_),
    .B1(_02723_),
    .C1(_02741_),
    .X(_02742_));
 sky130_fd_sc_hd__a211o_1 _08265_ (.A1(\_231_[21] ),
    .A2(_02730_),
    .B1(_02712_),
    .C1(_02742_),
    .X(_00328_));
 sky130_fd_sc_hd__or2_1 _08266_ (.A(\_164_[22] ),
    .B(_02736_),
    .X(_02743_));
 sky130_fd_sc_hd__o211a_1 _08267_ (.A1(\_228_[22] ),
    .A2(_02733_),
    .B1(_02723_),
    .C1(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__a211o_1 _08268_ (.A1(\_231_[22] ),
    .A2(_02730_),
    .B1(_02712_),
    .C1(_02744_),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _08269_ (.A0(\_164_[23] ),
    .A1(\_228_[23] ),
    .S(_02687_),
    .X(_02745_));
 sky130_fd_sc_hd__or2_1 _08270_ (.A(_02686_),
    .B(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__o211a_1 _08271_ (.A1(\_231_[23] ),
    .A2(_02706_),
    .B1(_02695_),
    .C1(_02746_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _08272_ (.A0(\_164_[24] ),
    .A1(\_228_[24] ),
    .S(_02687_),
    .X(_02747_));
 sky130_fd_sc_hd__or2_1 _08273_ (.A(_02686_),
    .B(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__o211a_1 _08274_ (.A1(\_231_[24] ),
    .A2(_02706_),
    .B1(_02695_),
    .C1(_02748_),
    .X(_00331_));
 sky130_fd_sc_hd__buf_2 _08275_ (.A(_01404_),
    .X(_02749_));
 sky130_fd_sc_hd__buf_4 _08276_ (.A(_01518_),
    .X(_02750_));
 sky130_fd_sc_hd__mux2_1 _08277_ (.A0(\_164_[25] ),
    .A1(\_228_[25] ),
    .S(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__or2_1 _08278_ (.A(_02749_),
    .B(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__o211a_1 _08279_ (.A1(\_231_[25] ),
    .A2(_02706_),
    .B1(_02695_),
    .C1(_02752_),
    .X(_00332_));
 sky130_fd_sc_hd__clkbuf_4 _08280_ (.A(_02711_),
    .X(_02753_));
 sky130_fd_sc_hd__or2_1 _08281_ (.A(\_164_[26] ),
    .B(_02736_),
    .X(_02754_));
 sky130_fd_sc_hd__o211a_1 _08282_ (.A1(\_228_[26] ),
    .A2(_02733_),
    .B1(_02723_),
    .C1(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__a211o_1 _08283_ (.A1(\_231_[26] ),
    .A2(_02730_),
    .B1(_02753_),
    .C1(_02755_),
    .X(_00333_));
 sky130_fd_sc_hd__or2_1 _08284_ (.A(\_164_[27] ),
    .B(_02736_),
    .X(_02756_));
 sky130_fd_sc_hd__o211a_1 _08285_ (.A1(\_228_[27] ),
    .A2(_02733_),
    .B1(_02723_),
    .C1(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__a211o_1 _08286_ (.A1(\_231_[27] ),
    .A2(_02730_),
    .B1(_02753_),
    .C1(_02757_),
    .X(_00334_));
 sky130_fd_sc_hd__or2_1 _08287_ (.A(\_164_[28] ),
    .B(_02736_),
    .X(_02758_));
 sky130_fd_sc_hd__o211a_1 _08288_ (.A1(\_228_[28] ),
    .A2(_02733_),
    .B1(_02723_),
    .C1(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__a211o_1 _08289_ (.A1(\_231_[28] ),
    .A2(_02730_),
    .B1(_02753_),
    .C1(_02759_),
    .X(_00335_));
 sky130_fd_sc_hd__buf_2 _08290_ (.A(_01420_),
    .X(_02760_));
 sky130_fd_sc_hd__or2_1 _08291_ (.A(\_164_[29] ),
    .B(_02736_),
    .X(_02761_));
 sky130_fd_sc_hd__o211a_1 _08292_ (.A1(\_228_[29] ),
    .A2(_02733_),
    .B1(_02760_),
    .C1(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__a211o_1 _08293_ (.A1(\_231_[29] ),
    .A2(_02730_),
    .B1(_02753_),
    .C1(_02762_),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _08294_ (.A0(\_164_[30] ),
    .A1(\_228_[30] ),
    .S(_02750_),
    .X(_02763_));
 sky130_fd_sc_hd__or2_1 _08295_ (.A(_02749_),
    .B(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__o211a_1 _08296_ (.A1(\_231_[30] ),
    .A2(_02706_),
    .B1(_02695_),
    .C1(_02764_),
    .X(_00337_));
 sky130_fd_sc_hd__clkbuf_4 _08297_ (.A(_01480_),
    .X(_02765_));
 sky130_fd_sc_hd__mux2_1 _08298_ (.A0(\_164_[31] ),
    .A1(\_228_[31] ),
    .S(_02750_),
    .X(_02766_));
 sky130_fd_sc_hd__or2_1 _08299_ (.A(_02749_),
    .B(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__o211a_1 _08300_ (.A1(\_231_[31] ),
    .A2(_02706_),
    .B1(_02765_),
    .C1(_02767_),
    .X(_00338_));
 sky130_fd_sc_hd__buf_4 _08301_ (.A(\_225_[0] ),
    .X(_02768_));
 sky130_fd_sc_hd__or2_1 _08302_ (.A(net36),
    .B(_02736_),
    .X(_02769_));
 sky130_fd_sc_hd__o211a_1 _08303_ (.A1(_02768_),
    .A2(_02733_),
    .B1(_02760_),
    .C1(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__a211o_1 _08304_ (.A1(\_228_[0] ),
    .A2(_02730_),
    .B1(_02753_),
    .C1(_02770_),
    .X(_00339_));
 sky130_fd_sc_hd__clkbuf_4 _08305_ (.A(_01799_),
    .X(_02771_));
 sky130_fd_sc_hd__buf_4 _08306_ (.A(\_225_[1] ),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _08307_ (.A0(net47),
    .A1(_02772_),
    .S(_02750_),
    .X(_02773_));
 sky130_fd_sc_hd__or2_1 _08308_ (.A(_02749_),
    .B(_02773_),
    .X(_02774_));
 sky130_fd_sc_hd__o211a_1 _08309_ (.A1(\_228_[1] ),
    .A2(_02771_),
    .B1(_02765_),
    .C1(_02774_),
    .X(_00340_));
 sky130_fd_sc_hd__buf_2 _08310_ (.A(_01406_),
    .X(_02775_));
 sky130_fd_sc_hd__buf_4 _08311_ (.A(\_225_[2] ),
    .X(_02776_));
 sky130_fd_sc_hd__or2_1 _08312_ (.A(net58),
    .B(_02736_),
    .X(_02777_));
 sky130_fd_sc_hd__o211a_1 _08313_ (.A1(_02776_),
    .A2(_02733_),
    .B1(_02760_),
    .C1(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__a211o_1 _08314_ (.A1(\_228_[2] ),
    .A2(_02775_),
    .B1(_02753_),
    .C1(_02778_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _08315_ (.A0(net61),
    .A1(\_225_[3] ),
    .S(_02750_),
    .X(_02779_));
 sky130_fd_sc_hd__or2_1 _08316_ (.A(_02749_),
    .B(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__o211a_1 _08317_ (.A1(\_228_[3] ),
    .A2(_02771_),
    .B1(_02765_),
    .C1(_02780_),
    .X(_00342_));
 sky130_fd_sc_hd__clkbuf_4 _08318_ (.A(\_225_[4] ),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _08319_ (.A0(net62),
    .A1(_02781_),
    .S(_02750_),
    .X(_02782_));
 sky130_fd_sc_hd__or2_1 _08320_ (.A(_02749_),
    .B(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__o211a_1 _08321_ (.A1(\_228_[4] ),
    .A2(_02771_),
    .B1(_02765_),
    .C1(_02783_),
    .X(_00343_));
 sky130_fd_sc_hd__clkbuf_4 _08322_ (.A(\_225_[5] ),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _08323_ (.A0(net63),
    .A1(_02784_),
    .S(_02750_),
    .X(_02785_));
 sky130_fd_sc_hd__or2_1 _08324_ (.A(_02749_),
    .B(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__o211a_1 _08325_ (.A1(\_228_[5] ),
    .A2(_02771_),
    .B1(_02765_),
    .C1(_02786_),
    .X(_00344_));
 sky130_fd_sc_hd__clkbuf_4 _08326_ (.A(\_225_[6] ),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _08327_ (.A0(net64),
    .A1(_02787_),
    .S(_02750_),
    .X(_02788_));
 sky130_fd_sc_hd__or2_1 _08328_ (.A(_02749_),
    .B(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__o211a_1 _08329_ (.A1(\_228_[6] ),
    .A2(_02771_),
    .B1(_02765_),
    .C1(_02789_),
    .X(_00345_));
 sky130_fd_sc_hd__clkbuf_4 _08330_ (.A(\_225_[7] ),
    .X(_02790_));
 sky130_fd_sc_hd__buf_2 _08331_ (.A(_01437_),
    .X(_02791_));
 sky130_fd_sc_hd__or2_1 _08332_ (.A(net65),
    .B(_02736_),
    .X(_02792_));
 sky130_fd_sc_hd__o211a_1 _08333_ (.A1(_02790_),
    .A2(_02791_),
    .B1(_02760_),
    .C1(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__a211o_1 _08334_ (.A1(\_228_[7] ),
    .A2(_02775_),
    .B1(_02753_),
    .C1(_02793_),
    .X(_00346_));
 sky130_fd_sc_hd__buf_4 _08335_ (.A(\_225_[8] ),
    .X(_02794_));
 sky130_fd_sc_hd__mux2_1 _08336_ (.A0(net66),
    .A1(_02794_),
    .S(_02750_),
    .X(_02795_));
 sky130_fd_sc_hd__or2_1 _08337_ (.A(_02749_),
    .B(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__o211a_1 _08338_ (.A1(\_228_[8] ),
    .A2(_02771_),
    .B1(_02765_),
    .C1(_02796_),
    .X(_00347_));
 sky130_fd_sc_hd__clkbuf_4 _08339_ (.A(\_225_[9] ),
    .X(_02797_));
 sky130_fd_sc_hd__clkbuf_2 _08340_ (.A(_01339_),
    .X(_02798_));
 sky130_fd_sc_hd__or2_1 _08341_ (.A(net67),
    .B(_02798_),
    .X(_02799_));
 sky130_fd_sc_hd__o211a_1 _08342_ (.A1(_02797_),
    .A2(_02791_),
    .B1(_02760_),
    .C1(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__a211o_1 _08343_ (.A1(\_228_[9] ),
    .A2(_02775_),
    .B1(_02753_),
    .C1(_02800_),
    .X(_00348_));
 sky130_fd_sc_hd__clkbuf_4 _08344_ (.A(\_225_[10] ),
    .X(_02801_));
 sky130_fd_sc_hd__or2_1 _08345_ (.A(net37),
    .B(_02798_),
    .X(_02802_));
 sky130_fd_sc_hd__o211a_1 _08346_ (.A1(_02801_),
    .A2(_02791_),
    .B1(_02760_),
    .C1(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__a211o_1 _08347_ (.A1(\_228_[10] ),
    .A2(_02775_),
    .B1(_02753_),
    .C1(_02803_),
    .X(_00349_));
 sky130_fd_sc_hd__clkbuf_4 _08348_ (.A(\_225_[11] ),
    .X(_02804_));
 sky130_fd_sc_hd__or2_1 _08349_ (.A(net38),
    .B(_02798_),
    .X(_02805_));
 sky130_fd_sc_hd__o211a_1 _08350_ (.A1(_02804_),
    .A2(_02791_),
    .B1(_02760_),
    .C1(_02805_),
    .X(_02806_));
 sky130_fd_sc_hd__a211o_1 _08351_ (.A1(\_228_[11] ),
    .A2(_02775_),
    .B1(_02753_),
    .C1(_02806_),
    .X(_00350_));
 sky130_fd_sc_hd__clkbuf_4 _08352_ (.A(\_225_[12] ),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _08353_ (.A0(net39),
    .A1(_02807_),
    .S(_02750_),
    .X(_02808_));
 sky130_fd_sc_hd__or2_1 _08354_ (.A(_02749_),
    .B(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__o211a_1 _08355_ (.A1(\_228_[12] ),
    .A2(_02771_),
    .B1(_02765_),
    .C1(_02809_),
    .X(_00351_));
 sky130_fd_sc_hd__clkbuf_4 _08356_ (.A(_02711_),
    .X(_02810_));
 sky130_fd_sc_hd__clkbuf_4 _08357_ (.A(\_225_[13] ),
    .X(_02811_));
 sky130_fd_sc_hd__or2_1 _08358_ (.A(net40),
    .B(_02798_),
    .X(_02812_));
 sky130_fd_sc_hd__o211a_1 _08359_ (.A1(_02811_),
    .A2(_02791_),
    .B1(_02760_),
    .C1(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__a211o_1 _08360_ (.A1(\_228_[13] ),
    .A2(_02775_),
    .B1(_02810_),
    .C1(_02813_),
    .X(_00352_));
 sky130_fd_sc_hd__clkbuf_4 _08361_ (.A(\_225_[14] ),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_1 _08362_ (.A0(net41),
    .A1(_02814_),
    .S(_01353_),
    .X(_02815_));
 sky130_fd_sc_hd__or2_1 _08363_ (.A(_02002_),
    .B(_02815_),
    .X(_02816_));
 sky130_fd_sc_hd__o211a_1 _08364_ (.A1(\_228_[14] ),
    .A2(_02771_),
    .B1(_02765_),
    .C1(_02816_),
    .X(_00353_));
 sky130_fd_sc_hd__buf_4 _08365_ (.A(\_225_[15] ),
    .X(_02817_));
 sky130_fd_sc_hd__or2_1 _08366_ (.A(net42),
    .B(_02798_),
    .X(_02818_));
 sky130_fd_sc_hd__o211a_1 _08367_ (.A1(_02817_),
    .A2(_02791_),
    .B1(_02760_),
    .C1(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__a211o_1 _08368_ (.A1(\_228_[15] ),
    .A2(_02775_),
    .B1(_02810_),
    .C1(_02819_),
    .X(_00354_));
 sky130_fd_sc_hd__clkbuf_4 _08369_ (.A(\_225_[16] ),
    .X(_02820_));
 sky130_fd_sc_hd__or2_1 _08370_ (.A(net43),
    .B(_02798_),
    .X(_02821_));
 sky130_fd_sc_hd__o211a_1 _08371_ (.A1(_02820_),
    .A2(_02791_),
    .B1(_02760_),
    .C1(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__a211o_1 _08372_ (.A1(\_228_[16] ),
    .A2(_02775_),
    .B1(_02810_),
    .C1(_02822_),
    .X(_00355_));
 sky130_fd_sc_hd__clkbuf_4 _08373_ (.A(\_225_[17] ),
    .X(_02823_));
 sky130_fd_sc_hd__clkbuf_4 _08374_ (.A(_01411_),
    .X(_02824_));
 sky130_fd_sc_hd__or2_1 _08375_ (.A(net44),
    .B(_02798_),
    .X(_02825_));
 sky130_fd_sc_hd__o211a_1 _08376_ (.A1(_02823_),
    .A2(_02791_),
    .B1(_02824_),
    .C1(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__a211o_1 _08377_ (.A1(\_228_[17] ),
    .A2(_02775_),
    .B1(_02810_),
    .C1(_02826_),
    .X(_00356_));
 sky130_fd_sc_hd__buf_4 _08378_ (.A(\_225_[18] ),
    .X(_02827_));
 sky130_fd_sc_hd__or2_1 _08379_ (.A(net45),
    .B(_02798_),
    .X(_02828_));
 sky130_fd_sc_hd__o211a_1 _08380_ (.A1(_02827_),
    .A2(_02791_),
    .B1(_02824_),
    .C1(_02828_),
    .X(_02829_));
 sky130_fd_sc_hd__a211o_1 _08381_ (.A1(\_228_[18] ),
    .A2(_02775_),
    .B1(_02810_),
    .C1(_02829_),
    .X(_00357_));
 sky130_fd_sc_hd__buf_4 _08382_ (.A(\_225_[19] ),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_1 _08383_ (.A0(net46),
    .A1(_02830_),
    .S(_01353_),
    .X(_02831_));
 sky130_fd_sc_hd__or2_1 _08384_ (.A(_02002_),
    .B(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__o211a_1 _08385_ (.A1(\_228_[19] ),
    .A2(_02771_),
    .B1(_02765_),
    .C1(_02832_),
    .X(_00358_));
 sky130_fd_sc_hd__buf_6 _08386_ (.A(_01423_),
    .X(_02833_));
 sky130_fd_sc_hd__clkbuf_4 _08387_ (.A(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__clkbuf_4 _08388_ (.A(\_225_[20] ),
    .X(_02835_));
 sky130_fd_sc_hd__mux2_1 _08389_ (.A0(net48),
    .A1(_02835_),
    .S(_01353_),
    .X(_02836_));
 sky130_fd_sc_hd__or2_1 _08390_ (.A(_02002_),
    .B(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__o211a_1 _08391_ (.A1(\_228_[20] ),
    .A2(_02771_),
    .B1(_02834_),
    .C1(_02837_),
    .X(_00359_));
 sky130_fd_sc_hd__clkbuf_4 _08392_ (.A(_01406_),
    .X(_02838_));
 sky130_fd_sc_hd__buf_4 _08393_ (.A(\_225_[21] ),
    .X(_02839_));
 sky130_fd_sc_hd__or2_1 _08394_ (.A(net49),
    .B(_02798_),
    .X(_02840_));
 sky130_fd_sc_hd__o211a_1 _08395_ (.A1(_02839_),
    .A2(_02791_),
    .B1(_02824_),
    .C1(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__a211o_1 _08396_ (.A1(\_228_[21] ),
    .A2(_02838_),
    .B1(_02810_),
    .C1(_02841_),
    .X(_00360_));
 sky130_fd_sc_hd__buf_4 _08397_ (.A(\_225_[22] ),
    .X(_02842_));
 sky130_fd_sc_hd__or2_1 _08398_ (.A(net50),
    .B(_02798_),
    .X(_02843_));
 sky130_fd_sc_hd__o211a_1 _08399_ (.A1(_02842_),
    .A2(_01801_),
    .B1(_02824_),
    .C1(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__a211o_1 _08400_ (.A1(\_228_[22] ),
    .A2(_02838_),
    .B1(_02810_),
    .C1(_02844_),
    .X(_00361_));
 sky130_fd_sc_hd__buf_4 _08401_ (.A(_01799_),
    .X(_02845_));
 sky130_fd_sc_hd__buf_6 _08402_ (.A(\_225_[23] ),
    .X(_02846_));
 sky130_fd_sc_hd__mux2_1 _08403_ (.A0(net51),
    .A1(_02846_),
    .S(_01353_),
    .X(_02847_));
 sky130_fd_sc_hd__or2_1 _08404_ (.A(_02002_),
    .B(_02847_),
    .X(_02848_));
 sky130_fd_sc_hd__o211a_1 _08405_ (.A1(\_228_[23] ),
    .A2(_02845_),
    .B1(_02834_),
    .C1(_02848_),
    .X(_00362_));
 sky130_fd_sc_hd__buf_4 _08406_ (.A(\_225_[24] ),
    .X(_02849_));
 sky130_fd_sc_hd__or2_1 _08407_ (.A(net52),
    .B(_01519_),
    .X(_02850_));
 sky130_fd_sc_hd__o211a_1 _08408_ (.A1(_02849_),
    .A2(_01801_),
    .B1(_02824_),
    .C1(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__a211o_1 _08409_ (.A1(\_228_[24] ),
    .A2(_02838_),
    .B1(_02810_),
    .C1(_02851_),
    .X(_00363_));
 sky130_fd_sc_hd__buf_4 _08410_ (.A(\_225_[25] ),
    .X(_02852_));
 sky130_fd_sc_hd__or2_1 _08411_ (.A(net53),
    .B(_01519_),
    .X(_02853_));
 sky130_fd_sc_hd__o211a_1 _08412_ (.A1(_02852_),
    .A2(_01801_),
    .B1(_02824_),
    .C1(_02853_),
    .X(_02854_));
 sky130_fd_sc_hd__a211o_1 _08413_ (.A1(\_228_[25] ),
    .A2(_02838_),
    .B1(_02810_),
    .C1(_02854_),
    .X(_00364_));
 sky130_fd_sc_hd__buf_6 _08414_ (.A(\_225_[26] ),
    .X(_02855_));
 sky130_fd_sc_hd__mux2_1 _08415_ (.A0(net54),
    .A1(_02855_),
    .S(_01353_),
    .X(_02856_));
 sky130_fd_sc_hd__or2_1 _08416_ (.A(_02002_),
    .B(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__o211a_1 _08417_ (.A1(\_228_[26] ),
    .A2(_02845_),
    .B1(_02834_),
    .C1(_02857_),
    .X(_00365_));
 sky130_fd_sc_hd__buf_6 _08418_ (.A(\_225_[27] ),
    .X(_02858_));
 sky130_fd_sc_hd__or2_1 _08419_ (.A(net55),
    .B(_01519_),
    .X(_02859_));
 sky130_fd_sc_hd__o211a_1 _08420_ (.A1(_02858_),
    .A2(_01801_),
    .B1(_02824_),
    .C1(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__a211o_1 _08421_ (.A1(\_228_[27] ),
    .A2(_02838_),
    .B1(_02810_),
    .C1(_02860_),
    .X(_00366_));
 sky130_fd_sc_hd__clkbuf_4 _08422_ (.A(_02711_),
    .X(_02861_));
 sky130_fd_sc_hd__buf_4 _08423_ (.A(\_225_[28] ),
    .X(_02862_));
 sky130_fd_sc_hd__or2_1 _08424_ (.A(net56),
    .B(_01519_),
    .X(_02863_));
 sky130_fd_sc_hd__o211a_1 _08425_ (.A1(_02862_),
    .A2(_01801_),
    .B1(_02824_),
    .C1(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__a211o_1 _08426_ (.A1(\_228_[28] ),
    .A2(_02838_),
    .B1(_02861_),
    .C1(_02864_),
    .X(_00367_));
 sky130_fd_sc_hd__buf_4 _08427_ (.A(\_225_[29] ),
    .X(_02865_));
 sky130_fd_sc_hd__or2_1 _08428_ (.A(net57),
    .B(_01519_),
    .X(_02866_));
 sky130_fd_sc_hd__o211a_1 _08429_ (.A1(_02865_),
    .A2(_01801_),
    .B1(_02824_),
    .C1(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__a211o_1 _08430_ (.A1(\_228_[29] ),
    .A2(_02838_),
    .B1(_02861_),
    .C1(_02867_),
    .X(_00368_));
 sky130_fd_sc_hd__buf_4 _08431_ (.A(\_225_[30] ),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _08432_ (.A0(net59),
    .A1(_02868_),
    .S(_01353_),
    .X(_02869_));
 sky130_fd_sc_hd__or2_1 _08433_ (.A(_02002_),
    .B(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__o211a_1 _08434_ (.A1(\_228_[30] ),
    .A2(_02845_),
    .B1(_02834_),
    .C1(_02870_),
    .X(_00369_));
 sky130_fd_sc_hd__buf_4 _08435_ (.A(\_225_[31] ),
    .X(_02871_));
 sky130_fd_sc_hd__or2_1 _08436_ (.A(net60),
    .B(_01519_),
    .X(_02872_));
 sky130_fd_sc_hd__o211a_1 _08437_ (.A1(_02871_),
    .A2(_01801_),
    .B1(_02824_),
    .C1(_02872_),
    .X(_02873_));
 sky130_fd_sc_hd__a211o_1 _08438_ (.A1(\_228_[31] ),
    .A2(_02838_),
    .B1(_02861_),
    .C1(_02873_),
    .X(_00370_));
 sky130_fd_sc_hd__xnor2_1 _08439_ (.A(_02811_),
    .B(_02776_),
    .Y(_02874_));
 sky130_fd_sc_hd__xnor2_2 _08440_ (.A(_02842_),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__xnor2_1 _08441_ (.A(\_185_[0] ),
    .B(_02875_),
    .Y(_02876_));
 sky130_fd_sc_hd__xnor2_1 _08442_ (.A(_01714_),
    .B(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__nand2_1 _08443_ (.A(_01719_),
    .B(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__or2_1 _08444_ (.A(_01719_),
    .B(_02877_),
    .X(_02879_));
 sky130_fd_sc_hd__nand2_1 _08445_ (.A(_02878_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__a21o_1 _08446_ (.A1(\_228_[0] ),
    .A2(\_231_[0] ),
    .B1(_02768_),
    .X(_02881_));
 sky130_fd_sc_hd__o21a_1 _08447_ (.A1(\_228_[0] ),
    .A2(\_231_[0] ),
    .B1(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__xnor2_1 _08448_ (.A(_02880_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__nand2_1 _08449_ (.A(\_170_[0] ),
    .B(_02768_),
    .Y(_02884_));
 sky130_fd_sc_hd__or2_1 _08450_ (.A(\_170_[0] ),
    .B(_02768_),
    .X(_02885_));
 sky130_fd_sc_hd__nand2_1 _08451_ (.A(_02884_),
    .B(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__nand2_1 _08452_ (.A(_02404_),
    .B(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__o211a_1 _08453_ (.A1(_02380_),
    .A2(_02883_),
    .B1(_02887_),
    .C1(_02202_),
    .X(_02888_));
 sky130_fd_sc_hd__a211o_1 _08454_ (.A1(_02768_),
    .A2(_02838_),
    .B1(_02861_),
    .C1(_02888_),
    .X(_00371_));
 sky130_fd_sc_hd__and2b_1 _08455_ (.A_N(_02880_),
    .B(_02882_),
    .X(_02889_));
 sky130_fd_sc_hd__inv_2 _08456_ (.A(_01727_),
    .Y(_02890_));
 sky130_fd_sc_hd__xnor2_1 _08457_ (.A(_02814_),
    .B(\_225_[3] ),
    .Y(_02891_));
 sky130_fd_sc_hd__xnor2_2 _08458_ (.A(_02846_),
    .B(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__xnor2_1 _08459_ (.A(\_185_[1] ),
    .B(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__xnor2_1 _08460_ (.A(_02890_),
    .B(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__inv_2 _08461_ (.A(_01714_),
    .Y(_02895_));
 sky130_fd_sc_hd__nand2_1 _08462_ (.A(\_185_[0] ),
    .B(_02875_),
    .Y(_02896_));
 sky130_fd_sc_hd__o21a_1 _08463_ (.A1(_02895_),
    .A2(_02876_),
    .B1(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__xor2_1 _08464_ (.A(_02894_),
    .B(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__xnor2_1 _08465_ (.A(_01734_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__xor2_1 _08466_ (.A(_02878_),
    .B(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__a21o_1 _08467_ (.A1(\_228_[1] ),
    .A2(\_231_[1] ),
    .B1(_02772_),
    .X(_02901_));
 sky130_fd_sc_hd__o21a_1 _08468_ (.A1(\_228_[1] ),
    .A2(\_231_[1] ),
    .B1(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__xor2_1 _08469_ (.A(_02900_),
    .B(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__and2_1 _08470_ (.A(_02889_),
    .B(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__o21ai_1 _08471_ (.A1(_02889_),
    .A2(_02903_),
    .B1(_01518_),
    .Y(_02905_));
 sky130_fd_sc_hd__xor2_2 _08472_ (.A(\_170_[1] ),
    .B(_02772_),
    .X(_02906_));
 sky130_fd_sc_hd__xnor2_1 _08473_ (.A(_02884_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__a2bb2o_1 _08474_ (.A1_N(_02904_),
    .A2_N(_02905_),
    .B1(_01269_),
    .B2(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_1 _08475_ (.A0(_02772_),
    .A1(_02908_),
    .S(_01411_),
    .X(_02909_));
 sky130_fd_sc_hd__or2_1 _08476_ (.A(_01710_),
    .B(_02909_),
    .X(_02910_));
 sky130_fd_sc_hd__clkbuf_1 _08477_ (.A(_02910_),
    .X(_00372_));
 sky130_fd_sc_hd__inv_2 _08478_ (.A(_01755_),
    .Y(_02911_));
 sky130_fd_sc_hd__xnor2_1 _08479_ (.A(_02817_),
    .B(_02781_),
    .Y(_02912_));
 sky130_fd_sc_hd__xnor2_1 _08480_ (.A(_02849_),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__xnor2_1 _08481_ (.A(\_185_[2] ),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__xnor2_1 _08482_ (.A(_02911_),
    .B(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__nand2_1 _08483_ (.A(\_185_[1] ),
    .B(_02892_),
    .Y(_02916_));
 sky130_fd_sc_hd__o21a_1 _08484_ (.A1(_02890_),
    .A2(_02893_),
    .B1(_02916_),
    .X(_02917_));
 sky130_fd_sc_hd__xor2_1 _08485_ (.A(_02915_),
    .B(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__xnor2_1 _08486_ (.A(_01762_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__nor2_1 _08487_ (.A(_02894_),
    .B(_02897_),
    .Y(_02920_));
 sky130_fd_sc_hd__a21oi_1 _08488_ (.A1(_01734_),
    .A2(_02898_),
    .B1(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__xnor2_1 _08489_ (.A(_02919_),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__a21o_1 _08490_ (.A1(\_228_[2] ),
    .A2(\_231_[2] ),
    .B1(_02776_),
    .X(_02923_));
 sky130_fd_sc_hd__o21a_1 _08491_ (.A1(\_228_[2] ),
    .A2(\_231_[2] ),
    .B1(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__xnor2_2 _08492_ (.A(_02922_),
    .B(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__nor2_1 _08493_ (.A(_02878_),
    .B(_02899_),
    .Y(_02926_));
 sky130_fd_sc_hd__a21o_1 _08494_ (.A1(_02900_),
    .A2(_02902_),
    .B1(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__xor2_2 _08495_ (.A(_02925_),
    .B(_02927_),
    .X(_02928_));
 sky130_fd_sc_hd__nand2_1 _08496_ (.A(_02904_),
    .B(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__o21a_1 _08497_ (.A1(_02904_),
    .A2(_02928_),
    .B1(_01302_),
    .X(_02930_));
 sky130_fd_sc_hd__and2_1 _08498_ (.A(\_170_[1] ),
    .B(_02772_),
    .X(_02931_));
 sky130_fd_sc_hd__a31oi_4 _08499_ (.A1(\_170_[0] ),
    .A2(_02768_),
    .A3(_02906_),
    .B1(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__and2_1 _08500_ (.A(\_170_[2] ),
    .B(_02776_),
    .X(_02933_));
 sky130_fd_sc_hd__nor2_1 _08501_ (.A(\_170_[2] ),
    .B(_02776_),
    .Y(_02934_));
 sky130_fd_sc_hd__nor2_1 _08502_ (.A(_02933_),
    .B(_02934_),
    .Y(_02935_));
 sky130_fd_sc_hd__xnor2_1 _08503_ (.A(_02932_),
    .B(_02935_),
    .Y(_02936_));
 sky130_fd_sc_hd__a22o_1 _08504_ (.A1(_02929_),
    .A2(_02930_),
    .B1(_02936_),
    .B2(_01269_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_1 _08505_ (.A0(_02776_),
    .A1(_02937_),
    .S(_01411_),
    .X(_02938_));
 sky130_fd_sc_hd__or2_1 _08506_ (.A(_01710_),
    .B(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__clkbuf_1 _08507_ (.A(_02939_),
    .X(_00373_));
 sky130_fd_sc_hd__or2_1 _08508_ (.A(\_170_[3] ),
    .B(\_225_[3] ),
    .X(_02940_));
 sky130_fd_sc_hd__nand2_1 _08509_ (.A(\_170_[3] ),
    .B(\_225_[3] ),
    .Y(_02941_));
 sky130_fd_sc_hd__nand2_1 _08510_ (.A(_02940_),
    .B(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__nand2_1 _08511_ (.A(\_170_[2] ),
    .B(_02776_),
    .Y(_02943_));
 sky130_fd_sc_hd__o21ai_1 _08512_ (.A1(_02932_),
    .A2(_02934_),
    .B1(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__xor2_1 _08513_ (.A(_02942_),
    .B(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__inv_2 _08514_ (.A(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__nor2_1 _08515_ (.A(_02919_),
    .B(_02921_),
    .Y(_02947_));
 sky130_fd_sc_hd__and2b_1 _08516_ (.A_N(_02922_),
    .B(_02924_),
    .X(_02948_));
 sky130_fd_sc_hd__inv_2 _08517_ (.A(_01781_),
    .Y(_02949_));
 sky130_fd_sc_hd__xnor2_1 _08518_ (.A(_02820_),
    .B(_02784_),
    .Y(_02950_));
 sky130_fd_sc_hd__xnor2_2 _08519_ (.A(_02852_),
    .B(_02950_),
    .Y(_02951_));
 sky130_fd_sc_hd__xnor2_1 _08520_ (.A(\_185_[3] ),
    .B(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__xnor2_1 _08521_ (.A(_02949_),
    .B(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__nand2_1 _08522_ (.A(\_185_[2] ),
    .B(_02913_),
    .Y(_02954_));
 sky130_fd_sc_hd__o21a_1 _08523_ (.A1(_02911_),
    .A2(_02914_),
    .B1(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__xor2_1 _08524_ (.A(_02953_),
    .B(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__xnor2_1 _08525_ (.A(_01789_),
    .B(_02956_),
    .Y(_02957_));
 sky130_fd_sc_hd__nor2_1 _08526_ (.A(_02915_),
    .B(_02917_),
    .Y(_02958_));
 sky130_fd_sc_hd__a21oi_1 _08527_ (.A1(_01762_),
    .A2(_02918_),
    .B1(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__xnor2_1 _08528_ (.A(_02957_),
    .B(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__a21o_1 _08529_ (.A1(\_228_[3] ),
    .A2(\_231_[3] ),
    .B1(\_225_[3] ),
    .X(_02961_));
 sky130_fd_sc_hd__o21a_1 _08530_ (.A1(\_228_[3] ),
    .A2(\_231_[3] ),
    .B1(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__xnor2_1 _08531_ (.A(_02960_),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__o21a_1 _08532_ (.A1(_02947_),
    .A2(_02948_),
    .B1(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__nor3_1 _08533_ (.A(_02947_),
    .B(_02948_),
    .C(_02963_),
    .Y(_02965_));
 sky130_fd_sc_hd__nand2_1 _08534_ (.A(_02925_),
    .B(_02927_),
    .Y(_02966_));
 sky130_fd_sc_hd__a21boi_1 _08535_ (.A1(_02904_),
    .A2(_02928_),
    .B1_N(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__o21a_1 _08536_ (.A1(_02964_),
    .A2(_02965_),
    .B1(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__nor3_1 _08537_ (.A(_02967_),
    .B(_02964_),
    .C(_02965_),
    .Y(_02969_));
 sky130_fd_sc_hd__nor3_1 _08538_ (.A(_01923_),
    .B(_02968_),
    .C(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__a211o_1 _08539_ (.A1(_01856_),
    .A2(_02946_),
    .B1(_02970_),
    .C1(_02355_),
    .X(_02971_));
 sky130_fd_sc_hd__o211a_1 _08540_ (.A1(\_225_[3] ),
    .A2(_02845_),
    .B1(_02834_),
    .C1(_02971_),
    .X(_00374_));
 sky130_fd_sc_hd__nor2_1 _08541_ (.A(\_170_[4] ),
    .B(_02781_),
    .Y(_02972_));
 sky130_fd_sc_hd__nand2_1 _08542_ (.A(\_170_[4] ),
    .B(_02781_),
    .Y(_02973_));
 sky130_fd_sc_hd__and2b_1 _08543_ (.A_N(_02972_),
    .B(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__o211ai_1 _08544_ (.A1(_02932_),
    .A2(_02934_),
    .B1(_02941_),
    .C1(_02943_),
    .Y(_02975_));
 sky130_fd_sc_hd__nand2_1 _08545_ (.A(_02940_),
    .B(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__xnor2_2 _08546_ (.A(_02974_),
    .B(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__nor2_1 _08547_ (.A(_02957_),
    .B(_02959_),
    .Y(_02978_));
 sky130_fd_sc_hd__and2b_1 _08548_ (.A_N(_02960_),
    .B(_02962_),
    .X(_02979_));
 sky130_fd_sc_hd__xnor2_1 _08549_ (.A(_02823_),
    .B(_02787_),
    .Y(_02980_));
 sky130_fd_sc_hd__xnor2_2 _08550_ (.A(_02855_),
    .B(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__xnor2_1 _08551_ (.A(\_185_[4] ),
    .B(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__xnor2_1 _08552_ (.A(_01835_),
    .B(_02982_),
    .Y(_02983_));
 sky130_fd_sc_hd__nand2_1 _08553_ (.A(\_185_[3] ),
    .B(_02951_),
    .Y(_02984_));
 sky130_fd_sc_hd__o21ai_1 _08554_ (.A1(_02949_),
    .A2(_02952_),
    .B1(_02984_),
    .Y(_02985_));
 sky130_fd_sc_hd__xnor2_1 _08555_ (.A(_02983_),
    .B(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hd__xnor2_1 _08556_ (.A(_01814_),
    .B(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__nor2_1 _08557_ (.A(_02953_),
    .B(_02955_),
    .Y(_02988_));
 sky130_fd_sc_hd__a21oi_1 _08558_ (.A1(_01789_),
    .A2(_02956_),
    .B1(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__xnor2_1 _08559_ (.A(_02987_),
    .B(_02989_),
    .Y(_02990_));
 sky130_fd_sc_hd__a21o_1 _08560_ (.A1(\_228_[4] ),
    .A2(\_231_[4] ),
    .B1(_02781_),
    .X(_02991_));
 sky130_fd_sc_hd__o21a_1 _08561_ (.A1(\_228_[4] ),
    .A2(\_231_[4] ),
    .B1(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__xnor2_1 _08562_ (.A(_02990_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__o21ai_1 _08563_ (.A1(_02978_),
    .A2(_02979_),
    .B1(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__or3_1 _08564_ (.A(_02978_),
    .B(_02979_),
    .C(_02993_),
    .X(_02995_));
 sky130_fd_sc_hd__and2_1 _08565_ (.A(_02994_),
    .B(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__nor2_1 _08566_ (.A(_02967_),
    .B(_02965_),
    .Y(_02997_));
 sky130_fd_sc_hd__o31a_1 _08567_ (.A1(_02964_),
    .A2(_02996_),
    .A3(_02997_),
    .B1(_01523_),
    .X(_02998_));
 sky130_fd_sc_hd__o21ai_1 _08568_ (.A1(_02964_),
    .A2(_02997_),
    .B1(_02996_),
    .Y(_02999_));
 sky130_fd_sc_hd__a221o_1 _08569_ (.A1(_02380_),
    .A2(_02977_),
    .B1(_02998_),
    .B2(_02999_),
    .C1(_01406_),
    .X(_03000_));
 sky130_fd_sc_hd__o211a_1 _08570_ (.A1(_02781_),
    .A2(_02845_),
    .B1(_02834_),
    .C1(_03000_),
    .X(_00375_));
 sky130_fd_sc_hd__nand2_1 _08571_ (.A(_02994_),
    .B(_02999_),
    .Y(_03001_));
 sky130_fd_sc_hd__nor2_1 _08572_ (.A(_02987_),
    .B(_02989_),
    .Y(_03002_));
 sky130_fd_sc_hd__and2b_1 _08573_ (.A_N(_02990_),
    .B(_02992_),
    .X(_03003_));
 sky130_fd_sc_hd__clkinv_2 _08574_ (.A(_01838_),
    .Y(_03004_));
 sky130_fd_sc_hd__xnor2_2 _08575_ (.A(_02827_),
    .B(_02790_),
    .Y(_03005_));
 sky130_fd_sc_hd__xnor2_4 _08576_ (.A(_02858_),
    .B(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__xnor2_4 _08577_ (.A(\_185_[5] ),
    .B(_03006_),
    .Y(_03007_));
 sky130_fd_sc_hd__xnor2_4 _08578_ (.A(_03004_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__nand2_1 _08579_ (.A(\_185_[4] ),
    .B(_02981_),
    .Y(_03009_));
 sky130_fd_sc_hd__o21a_1 _08580_ (.A1(_01835_),
    .A2(_02982_),
    .B1(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__xor2_4 _08581_ (.A(_03008_),
    .B(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__xnor2_2 _08582_ (.A(_01847_),
    .B(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__and2b_1 _08583_ (.A_N(_02983_),
    .B(_02985_),
    .X(_03013_));
 sky130_fd_sc_hd__a21oi_2 _08584_ (.A1(_01814_),
    .A2(_02986_),
    .B1(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__xnor2_2 _08585_ (.A(_03012_),
    .B(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__nor2_1 _08586_ (.A(\_228_[5] ),
    .B(\_231_[5] ),
    .Y(_03016_));
 sky130_fd_sc_hd__a21oi_2 _08587_ (.A1(\_228_[5] ),
    .A2(\_231_[5] ),
    .B1(_02784_),
    .Y(_03017_));
 sky130_fd_sc_hd__nor2_1 _08588_ (.A(_03016_),
    .B(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__xnor2_1 _08589_ (.A(_03015_),
    .B(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__nor3_1 _08590_ (.A(_03002_),
    .B(_03003_),
    .C(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__o21ai_1 _08591_ (.A1(_03002_),
    .A2(_03003_),
    .B1(_03019_),
    .Y(_03021_));
 sky130_fd_sc_hd__or2b_1 _08592_ (.A(_03020_),
    .B_N(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__and2_1 _08593_ (.A(_03001_),
    .B(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__o21ai_1 _08594_ (.A1(_03001_),
    .A2(_03022_),
    .B1(_01354_),
    .Y(_03024_));
 sky130_fd_sc_hd__or2_1 _08595_ (.A(\_170_[5] ),
    .B(_02784_),
    .X(_03025_));
 sky130_fd_sc_hd__nand2_1 _08596_ (.A(\_170_[5] ),
    .B(_02784_),
    .Y(_03026_));
 sky130_fd_sc_hd__nand2_1 _08597_ (.A(_03025_),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__o21a_1 _08598_ (.A1(_02972_),
    .A2(_02976_),
    .B1(_02973_),
    .X(_03028_));
 sky130_fd_sc_hd__xnor2_1 _08599_ (.A(_03027_),
    .B(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hd__inv_2 _08600_ (.A(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__o221a_1 _08601_ (.A1(_03023_),
    .A2(_03024_),
    .B1(_03030_),
    .B2(_01520_),
    .C1(_01439_),
    .X(_03031_));
 sky130_fd_sc_hd__a211o_1 _08602_ (.A1(_02784_),
    .A2(_02838_),
    .B1(_02861_),
    .C1(_03031_),
    .X(_00376_));
 sky130_fd_sc_hd__clkbuf_4 _08603_ (.A(_01406_),
    .X(_03032_));
 sky130_fd_sc_hd__inv_2 _08604_ (.A(_01867_),
    .Y(_03033_));
 sky130_fd_sc_hd__xnor2_1 _08605_ (.A(_02830_),
    .B(_02794_),
    .Y(_03034_));
 sky130_fd_sc_hd__xnor2_2 _08606_ (.A(_02862_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__xnor2_1 _08607_ (.A(\_185_[6] ),
    .B(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__xnor2_2 _08608_ (.A(_03033_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__nand2_1 _08609_ (.A(\_185_[5] ),
    .B(_03006_),
    .Y(_03038_));
 sky130_fd_sc_hd__o21ai_2 _08610_ (.A1(_03004_),
    .A2(_03007_),
    .B1(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__xnor2_4 _08611_ (.A(_03037_),
    .B(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__xnor2_4 _08612_ (.A(_01875_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__nor2_1 _08613_ (.A(_03008_),
    .B(_03010_),
    .Y(_03042_));
 sky130_fd_sc_hd__a21oi_4 _08614_ (.A1(_01847_),
    .A2(_03011_),
    .B1(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__xnor2_2 _08615_ (.A(_03041_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__nor2_1 _08616_ (.A(\_228_[6] ),
    .B(\_231_[6] ),
    .Y(_03045_));
 sky130_fd_sc_hd__a21oi_2 _08617_ (.A1(\_228_[6] ),
    .A2(\_231_[6] ),
    .B1(_02787_),
    .Y(_03046_));
 sky130_fd_sc_hd__nor2_1 _08618_ (.A(_03045_),
    .B(_03046_),
    .Y(_03047_));
 sky130_fd_sc_hd__xnor2_2 _08619_ (.A(_03044_),
    .B(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__o32ai_4 _08620_ (.A1(_03015_),
    .A2(_03016_),
    .A3(_03017_),
    .B1(_03014_),
    .B2(_03012_),
    .Y(_03049_));
 sky130_fd_sc_hd__xor2_2 _08621_ (.A(_03048_),
    .B(_03049_),
    .X(_03050_));
 sky130_fd_sc_hd__a21o_1 _08622_ (.A1(_02994_),
    .A2(_03021_),
    .B1(_03020_),
    .X(_03051_));
 sky130_fd_sc_hd__o21ai_1 _08623_ (.A1(_02999_),
    .A2(_03020_),
    .B1(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__xor2_1 _08624_ (.A(_03050_),
    .B(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__or2_1 _08625_ (.A(\_170_[6] ),
    .B(_02787_),
    .X(_03054_));
 sky130_fd_sc_hd__nand2_1 _08626_ (.A(\_170_[6] ),
    .B(_02787_),
    .Y(_03055_));
 sky130_fd_sc_hd__nand2_1 _08627_ (.A(_03054_),
    .B(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__nand2_1 _08628_ (.A(_02973_),
    .B(_03026_),
    .Y(_03057_));
 sky130_fd_sc_hd__a31o_1 _08629_ (.A1(_02940_),
    .A2(_02974_),
    .A3(_02975_),
    .B1(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__nand2_1 _08630_ (.A(_03025_),
    .B(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__xnor2_1 _08631_ (.A(_03056_),
    .B(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__nand2_1 _08632_ (.A(_02404_),
    .B(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__o211a_1 _08633_ (.A1(_02380_),
    .A2(_03053_),
    .B1(_03061_),
    .C1(_02202_),
    .X(_03062_));
 sky130_fd_sc_hd__a211o_1 _08634_ (.A1(_02787_),
    .A2(_03032_),
    .B1(_02861_),
    .C1(_03062_),
    .X(_00377_));
 sky130_fd_sc_hd__nor2_1 _08635_ (.A(\_170_[7] ),
    .B(_02790_),
    .Y(_03063_));
 sky130_fd_sc_hd__and2_1 _08636_ (.A(\_170_[7] ),
    .B(_02790_),
    .X(_03064_));
 sky130_fd_sc_hd__nor2_1 _08637_ (.A(_03063_),
    .B(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__and2_1 _08638_ (.A(\_170_[6] ),
    .B(_02787_),
    .X(_03066_));
 sky130_fd_sc_hd__a31o_1 _08639_ (.A1(_03025_),
    .A2(_03054_),
    .A3(_03058_),
    .B1(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__xnor2_1 _08640_ (.A(_03065_),
    .B(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__inv_2 _08641_ (.A(_03068_),
    .Y(_03069_));
 sky130_fd_sc_hd__o32ai_4 _08642_ (.A1(_03044_),
    .A2(_03045_),
    .A3(_03046_),
    .B1(_03043_),
    .B2(_03041_),
    .Y(_03070_));
 sky130_fd_sc_hd__xnor2_1 _08643_ (.A(_02835_),
    .B(_02797_),
    .Y(_03071_));
 sky130_fd_sc_hd__xnor2_2 _08644_ (.A(_02865_),
    .B(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hd__xnor2_1 _08645_ (.A(\_185_[7] ),
    .B(_03072_),
    .Y(_03073_));
 sky130_fd_sc_hd__xnor2_1 _08646_ (.A(_01927_),
    .B(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_1 _08647_ (.A(\_185_[6] ),
    .B(_03035_),
    .Y(_03075_));
 sky130_fd_sc_hd__o21a_1 _08648_ (.A1(_03033_),
    .A2(_03036_),
    .B1(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__xnor2_1 _08649_ (.A(_03074_),
    .B(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__xor2_2 _08650_ (.A(_01906_),
    .B(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__and2b_1 _08651_ (.A_N(_03037_),
    .B(_03039_),
    .X(_03079_));
 sky130_fd_sc_hd__a21oi_2 _08652_ (.A1(_01875_),
    .A2(_03040_),
    .B1(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__xnor2_2 _08653_ (.A(_03078_),
    .B(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__nor2_1 _08654_ (.A(\_228_[7] ),
    .B(\_231_[7] ),
    .Y(_03082_));
 sky130_fd_sc_hd__a21oi_1 _08655_ (.A1(\_228_[7] ),
    .A2(\_231_[7] ),
    .B1(_02790_),
    .Y(_03083_));
 sky130_fd_sc_hd__nor2_1 _08656_ (.A(_03082_),
    .B(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__xnor2_2 _08657_ (.A(_03081_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__xor2_2 _08658_ (.A(_03070_),
    .B(_03085_),
    .X(_03086_));
 sky130_fd_sc_hd__nand2_1 _08659_ (.A(_03048_),
    .B(_03049_),
    .Y(_03087_));
 sky130_fd_sc_hd__a21bo_1 _08660_ (.A1(_03050_),
    .A2(_03052_),
    .B1_N(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__xnor2_1 _08661_ (.A(_03086_),
    .B(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__nor2_1 _08662_ (.A(_01923_),
    .B(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__a211o_1 _08663_ (.A1(_01856_),
    .A2(_03069_),
    .B1(_03090_),
    .C1(_02355_),
    .X(_03091_));
 sky130_fd_sc_hd__o211a_1 _08664_ (.A1(_02790_),
    .A2(_02845_),
    .B1(_02834_),
    .C1(_03091_),
    .X(_00378_));
 sky130_fd_sc_hd__a21oi_1 _08665_ (.A1(_02904_),
    .A2(_02928_),
    .B1(_02964_),
    .Y(_03092_));
 sky130_fd_sc_hd__nand4b_1 _08666_ (.A_N(_03020_),
    .B(_03021_),
    .C(_03050_),
    .D(_03086_),
    .Y(_03093_));
 sky130_fd_sc_hd__nand2_1 _08667_ (.A(_02994_),
    .B(_02995_),
    .Y(_03094_));
 sky130_fd_sc_hd__a2111o_1 _08668_ (.A1(_02966_),
    .A2(_03092_),
    .B1(_03093_),
    .C1(_02965_),
    .D1(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__nor2_1 _08669_ (.A(_03070_),
    .B(_03085_),
    .Y(_03096_));
 sky130_fd_sc_hd__nand2_1 _08670_ (.A(_03050_),
    .B(_03086_),
    .Y(_03097_));
 sky130_fd_sc_hd__nand2_1 _08671_ (.A(_03070_),
    .B(_03085_),
    .Y(_03098_));
 sky130_fd_sc_hd__o221a_1 _08672_ (.A1(_03087_),
    .A2(_03096_),
    .B1(_03097_),
    .B2(_03051_),
    .C1(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__and2_1 _08673_ (.A(_03095_),
    .B(_03099_),
    .X(_03100_));
 sky130_fd_sc_hd__clkinv_2 _08674_ (.A(_01930_),
    .Y(_03101_));
 sky130_fd_sc_hd__xnor2_2 _08675_ (.A(_02839_),
    .B(_02801_),
    .Y(_03102_));
 sky130_fd_sc_hd__xnor2_4 _08676_ (.A(_02868_),
    .B(_03102_),
    .Y(_03103_));
 sky130_fd_sc_hd__xnor2_2 _08677_ (.A(\_185_[8] ),
    .B(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__xnor2_4 _08678_ (.A(_03101_),
    .B(_03104_),
    .Y(_03105_));
 sky130_fd_sc_hd__nand2_1 _08679_ (.A(\_185_[7] ),
    .B(_03072_),
    .Y(_03106_));
 sky130_fd_sc_hd__o21a_1 _08680_ (.A1(_01927_),
    .A2(_03073_),
    .B1(_03106_),
    .X(_03107_));
 sky130_fd_sc_hd__xor2_4 _08681_ (.A(_03105_),
    .B(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__xnor2_4 _08682_ (.A(_01939_),
    .B(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__o32a_2 _08683_ (.A1(_01904_),
    .A2(_01905_),
    .A3(_03077_),
    .B1(_03076_),
    .B2(_03074_),
    .X(_03110_));
 sky130_fd_sc_hd__xnor2_2 _08684_ (.A(_03109_),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__nor2_1 _08685_ (.A(\_228_[8] ),
    .B(\_231_[8] ),
    .Y(_03112_));
 sky130_fd_sc_hd__a21oi_2 _08686_ (.A1(\_228_[8] ),
    .A2(\_231_[8] ),
    .B1(_02794_),
    .Y(_03113_));
 sky130_fd_sc_hd__nor2_1 _08687_ (.A(_03112_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__xnor2_1 _08688_ (.A(_03111_),
    .B(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__o32a_1 _08689_ (.A1(_03081_),
    .A2(_03082_),
    .A3(_03083_),
    .B1(_03080_),
    .B2(_03078_),
    .X(_03116_));
 sky130_fd_sc_hd__xnor2_1 _08690_ (.A(_03115_),
    .B(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__xnor2_1 _08691_ (.A(_03100_),
    .B(_03117_),
    .Y(_03118_));
 sky130_fd_sc_hd__nor2_1 _08692_ (.A(\_170_[8] ),
    .B(_02794_),
    .Y(_03119_));
 sky130_fd_sc_hd__and2_1 _08693_ (.A(\_170_[8] ),
    .B(_02794_),
    .X(_03120_));
 sky130_fd_sc_hd__nor2_1 _08694_ (.A(_03119_),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__or2_1 _08695_ (.A(\_170_[7] ),
    .B(_02790_),
    .X(_03122_));
 sky130_fd_sc_hd__a311o_1 _08696_ (.A1(_03025_),
    .A2(_03054_),
    .A3(_03058_),
    .B1(_03064_),
    .C1(_03066_),
    .X(_03123_));
 sky130_fd_sc_hd__nand2_1 _08697_ (.A(_03122_),
    .B(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__xor2_1 _08698_ (.A(_03121_),
    .B(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__nor2_1 _08699_ (.A(_01778_),
    .B(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__a211o_1 _08700_ (.A1(_01355_),
    .A2(_03118_),
    .B1(_03126_),
    .C1(_02355_),
    .X(_03127_));
 sky130_fd_sc_hd__o211a_1 _08701_ (.A1(_02794_),
    .A2(_02845_),
    .B1(_02834_),
    .C1(_03127_),
    .X(_00379_));
 sky130_fd_sc_hd__or2_1 _08702_ (.A(\_170_[9] ),
    .B(_02797_),
    .X(_03128_));
 sky130_fd_sc_hd__nand2_1 _08703_ (.A(\_170_[9] ),
    .B(_02797_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand2_1 _08704_ (.A(_03128_),
    .B(_03129_),
    .Y(_03130_));
 sky130_fd_sc_hd__a31oi_2 _08705_ (.A1(_03122_),
    .A2(_03121_),
    .A3(_03123_),
    .B1(_03120_),
    .Y(_03131_));
 sky130_fd_sc_hd__xnor2_1 _08706_ (.A(_03130_),
    .B(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__inv_2 _08707_ (.A(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__or2b_1 _08708_ (.A(_03116_),
    .B_N(_03115_),
    .X(_03134_));
 sky130_fd_sc_hd__or2b_1 _08709_ (.A(_03100_),
    .B_N(_03117_),
    .X(_03135_));
 sky130_fd_sc_hd__o32ai_4 _08710_ (.A1(_03111_),
    .A2(_03112_),
    .A3(_03113_),
    .B1(_03110_),
    .B2(_03109_),
    .Y(_03136_));
 sky130_fd_sc_hd__xnor2_1 _08711_ (.A(_02842_),
    .B(_02804_),
    .Y(_03137_));
 sky130_fd_sc_hd__xnor2_2 _08712_ (.A(_02871_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__xnor2_1 _08713_ (.A(\_185_[9] ),
    .B(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__xnor2_1 _08714_ (.A(_01974_),
    .B(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__nand2_1 _08715_ (.A(\_185_[8] ),
    .B(_03103_),
    .Y(_03141_));
 sky130_fd_sc_hd__o21ai_1 _08716_ (.A1(_03101_),
    .A2(_03104_),
    .B1(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__xnor2_1 _08717_ (.A(_03140_),
    .B(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__xnor2_2 _08718_ (.A(_01960_),
    .B(_03143_),
    .Y(_03144_));
 sky130_fd_sc_hd__nor2_1 _08719_ (.A(_03105_),
    .B(_03107_),
    .Y(_03145_));
 sky130_fd_sc_hd__a21oi_2 _08720_ (.A1(_01939_),
    .A2(_03108_),
    .B1(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__xnor2_1 _08721_ (.A(_03144_),
    .B(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__nor2_1 _08722_ (.A(\_228_[9] ),
    .B(\_231_[9] ),
    .Y(_03148_));
 sky130_fd_sc_hd__a21oi_2 _08723_ (.A1(\_228_[9] ),
    .A2(\_231_[9] ),
    .B1(_02797_),
    .Y(_03149_));
 sky130_fd_sc_hd__nor2_1 _08724_ (.A(_03148_),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__xnor2_1 _08725_ (.A(_03147_),
    .B(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__xor2_1 _08726_ (.A(_03136_),
    .B(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__and3_1 _08727_ (.A(_03134_),
    .B(_03135_),
    .C(_03152_),
    .X(_03153_));
 sky130_fd_sc_hd__a21oi_1 _08728_ (.A1(_03134_),
    .A2(_03135_),
    .B1(_03152_),
    .Y(_03154_));
 sky130_fd_sc_hd__or3_1 _08729_ (.A(_01408_),
    .B(_03153_),
    .C(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__o211a_1 _08730_ (.A1(_01520_),
    .A2(_03133_),
    .B1(_03155_),
    .C1(_02202_),
    .X(_03156_));
 sky130_fd_sc_hd__a211o_1 _08731_ (.A1(_02797_),
    .A2(_03032_),
    .B1(_02861_),
    .C1(_03156_),
    .X(_00380_));
 sky130_fd_sc_hd__xnor2_1 _08732_ (.A(_02807_),
    .B(_02768_),
    .Y(_03157_));
 sky130_fd_sc_hd__xnor2_2 _08733_ (.A(_02846_),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__xnor2_1 _08734_ (.A(\_185_[10] ),
    .B(_03158_),
    .Y(_03159_));
 sky130_fd_sc_hd__xnor2_1 _08735_ (.A(_02006_),
    .B(_03159_),
    .Y(_03160_));
 sky130_fd_sc_hd__nand2_1 _08736_ (.A(\_185_[9] ),
    .B(_03138_),
    .Y(_03161_));
 sky130_fd_sc_hd__o21a_1 _08737_ (.A1(_01974_),
    .A2(_03139_),
    .B1(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__xor2_1 _08738_ (.A(_03160_),
    .B(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__xnor2_1 _08739_ (.A(_01985_),
    .B(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__and2b_1 _08740_ (.A_N(_03140_),
    .B(_03142_),
    .X(_03165_));
 sky130_fd_sc_hd__a21oi_1 _08741_ (.A1(_01960_),
    .A2(_03143_),
    .B1(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__xnor2_1 _08742_ (.A(_03164_),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__a21o_1 _08743_ (.A1(\_228_[10] ),
    .A2(\_231_[10] ),
    .B1(_02801_),
    .X(_03168_));
 sky130_fd_sc_hd__o21a_1 _08744_ (.A1(\_228_[10] ),
    .A2(\_231_[10] ),
    .B1(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__xnor2_1 _08745_ (.A(_03167_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__o32ai_2 _08746_ (.A1(_03147_),
    .A2(_03148_),
    .A3(_03149_),
    .B1(_03146_),
    .B2(_03144_),
    .Y(_03171_));
 sky130_fd_sc_hd__xor2_1 _08747_ (.A(_03170_),
    .B(_03171_),
    .X(_03172_));
 sky130_fd_sc_hd__nand2_1 _08748_ (.A(_03117_),
    .B(_03152_),
    .Y(_03173_));
 sky130_fd_sc_hd__nand2_1 _08749_ (.A(_03136_),
    .B(_03151_),
    .Y(_03174_));
 sky130_fd_sc_hd__nor2_1 _08750_ (.A(_03136_),
    .B(_03151_),
    .Y(_03175_));
 sky130_fd_sc_hd__a21o_1 _08751_ (.A1(_03134_),
    .A2(_03174_),
    .B1(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__o21ai_1 _08752_ (.A1(_03100_),
    .A2(_03173_),
    .B1(_03176_),
    .Y(_03177_));
 sky130_fd_sc_hd__xor2_1 _08753_ (.A(_03172_),
    .B(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__and2_1 _08754_ (.A(\_170_[10] ),
    .B(_02801_),
    .X(_03179_));
 sky130_fd_sc_hd__nor2_1 _08755_ (.A(\_170_[10] ),
    .B(_02801_),
    .Y(_03180_));
 sky130_fd_sc_hd__or2_1 _08756_ (.A(_03179_),
    .B(_03180_),
    .X(_03181_));
 sky130_fd_sc_hd__inv_2 _08757_ (.A(_03128_),
    .Y(_03182_));
 sky130_fd_sc_hd__a21oi_1 _08758_ (.A1(_03129_),
    .A2(_03131_),
    .B1(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__xor2_2 _08759_ (.A(_03181_),
    .B(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__nand2_1 _08760_ (.A(_02404_),
    .B(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__o211a_1 _08761_ (.A1(_02380_),
    .A2(_03178_),
    .B1(_03185_),
    .C1(_02202_),
    .X(_03186_));
 sky130_fd_sc_hd__a211o_1 _08762_ (.A1(_02801_),
    .A2(_03032_),
    .B1(_02861_),
    .C1(_03186_),
    .X(_00381_));
 sky130_fd_sc_hd__nand2_1 _08763_ (.A(_03170_),
    .B(_03171_),
    .Y(_03187_));
 sky130_fd_sc_hd__nand2_1 _08764_ (.A(_03172_),
    .B(_03177_),
    .Y(_03188_));
 sky130_fd_sc_hd__nor2_1 _08765_ (.A(_03164_),
    .B(_03166_),
    .Y(_03189_));
 sky130_fd_sc_hd__and2b_1 _08766_ (.A_N(_03167_),
    .B(_03169_),
    .X(_03190_));
 sky130_fd_sc_hd__xnor2_1 _08767_ (.A(_02811_),
    .B(_02772_),
    .Y(_03191_));
 sky130_fd_sc_hd__xnor2_2 _08768_ (.A(_02849_),
    .B(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__xnor2_1 _08769_ (.A(\_185_[11] ),
    .B(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__xnor2_1 _08770_ (.A(_02037_),
    .B(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__nand2_1 _08771_ (.A(\_185_[10] ),
    .B(_03158_),
    .Y(_03195_));
 sky130_fd_sc_hd__o21a_1 _08772_ (.A1(_02006_),
    .A2(_03159_),
    .B1(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__xnor2_1 _08773_ (.A(_03194_),
    .B(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__xor2_1 _08774_ (.A(_02017_),
    .B(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__nor2_1 _08775_ (.A(_03160_),
    .B(_03162_),
    .Y(_03199_));
 sky130_fd_sc_hd__a21oi_2 _08776_ (.A1(_01985_),
    .A2(_03163_),
    .B1(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__xnor2_1 _08777_ (.A(_03198_),
    .B(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hd__a21o_1 _08778_ (.A1(\_228_[11] ),
    .A2(\_231_[11] ),
    .B1(_02804_),
    .X(_03202_));
 sky130_fd_sc_hd__o21a_1 _08779_ (.A1(\_228_[11] ),
    .A2(\_231_[11] ),
    .B1(_03202_),
    .X(_03203_));
 sky130_fd_sc_hd__xnor2_1 _08780_ (.A(_03201_),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__nor3_1 _08781_ (.A(_03189_),
    .B(_03190_),
    .C(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__o21ai_1 _08782_ (.A1(_03189_),
    .A2(_03190_),
    .B1(_03204_),
    .Y(_03206_));
 sky130_fd_sc_hd__or2b_1 _08783_ (.A(_03205_),
    .B_N(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__a21oi_1 _08784_ (.A1(_03187_),
    .A2(_03188_),
    .B1(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__a31o_1 _08785_ (.A1(_03187_),
    .A2(_03188_),
    .A3(_03207_),
    .B1(_01923_),
    .X(_03209_));
 sky130_fd_sc_hd__and2_1 _08786_ (.A(\_170_[11] ),
    .B(_02804_),
    .X(_03210_));
 sky130_fd_sc_hd__nor2_1 _08787_ (.A(\_170_[11] ),
    .B(_02804_),
    .Y(_03211_));
 sky130_fd_sc_hd__or2_1 _08788_ (.A(_03210_),
    .B(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__a211oi_1 _08789_ (.A1(_03129_),
    .A2(_03131_),
    .B1(_03181_),
    .C1(_03182_),
    .Y(_03213_));
 sky130_fd_sc_hd__nor2_1 _08790_ (.A(_03179_),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__xnor2_2 _08791_ (.A(_03212_),
    .B(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__o21a_1 _08792_ (.A1(_01778_),
    .A2(_03215_),
    .B1(_01412_),
    .X(_03216_));
 sky130_fd_sc_hd__o21ai_1 _08793_ (.A1(_03208_),
    .A2(_03209_),
    .B1(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__o211a_1 _08794_ (.A1(_02804_),
    .A2(_02845_),
    .B1(_02834_),
    .C1(_03217_),
    .X(_00382_));
 sky130_fd_sc_hd__nor2_1 _08795_ (.A(_03194_),
    .B(_03196_),
    .Y(_03218_));
 sky130_fd_sc_hd__and2b_1 _08796_ (.A_N(_03197_),
    .B(_02017_),
    .X(_03219_));
 sky130_fd_sc_hd__xnor2_1 _08797_ (.A(_02814_),
    .B(_02776_),
    .Y(_03220_));
 sky130_fd_sc_hd__xnor2_2 _08798_ (.A(_02852_),
    .B(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__xnor2_1 _08799_ (.A(\_185_[12] ),
    .B(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__xnor2_1 _08800_ (.A(_02071_),
    .B(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__nand2_1 _08801_ (.A(\_185_[11] ),
    .B(_03192_),
    .Y(_03224_));
 sky130_fd_sc_hd__o21a_1 _08802_ (.A1(_02037_),
    .A2(_03193_),
    .B1(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__xor2_1 _08803_ (.A(_03223_),
    .B(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__xnor2_1 _08804_ (.A(_02048_),
    .B(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__o21ba_1 _08805_ (.A1(_03218_),
    .A2(_03219_),
    .B1_N(_03227_),
    .X(_03228_));
 sky130_fd_sc_hd__or3b_1 _08806_ (.A(_03218_),
    .B(_03219_),
    .C_N(_03227_),
    .X(_03229_));
 sky130_fd_sc_hd__or2b_1 _08807_ (.A(_03228_),
    .B_N(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__a21o_1 _08808_ (.A1(\_228_[12] ),
    .A2(\_231_[12] ),
    .B1(_02807_),
    .X(_03231_));
 sky130_fd_sc_hd__o21a_1 _08809_ (.A1(\_228_[12] ),
    .A2(\_231_[12] ),
    .B1(_03231_),
    .X(_03232_));
 sky130_fd_sc_hd__xnor2_1 _08810_ (.A(_03230_),
    .B(_03232_),
    .Y(_03233_));
 sky130_fd_sc_hd__or2b_1 _08811_ (.A(_03201_),
    .B_N(_03203_),
    .X(_03234_));
 sky130_fd_sc_hd__o21ai_1 _08812_ (.A1(_03198_),
    .A2(_03200_),
    .B1(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__xor2_1 _08813_ (.A(_03233_),
    .B(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__nand3b_1 _08814_ (.A_N(_03205_),
    .B(_03206_),
    .C(_03172_),
    .Y(_03237_));
 sky130_fd_sc_hd__or2_1 _08815_ (.A(_03173_),
    .B(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__o221a_1 _08816_ (.A1(_03187_),
    .A2(_03205_),
    .B1(_03237_),
    .B2(_03176_),
    .C1(_03206_),
    .X(_03239_));
 sky130_fd_sc_hd__o21ai_1 _08817_ (.A1(_03100_),
    .A2(_03238_),
    .B1(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__nand2_1 _08818_ (.A(_03236_),
    .B(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__or2_1 _08819_ (.A(_03236_),
    .B(_03240_),
    .X(_03242_));
 sky130_fd_sc_hd__or2_1 _08820_ (.A(\_170_[12] ),
    .B(_02807_),
    .X(_03243_));
 sky130_fd_sc_hd__nand2_1 _08821_ (.A(\_170_[12] ),
    .B(_02807_),
    .Y(_03244_));
 sky130_fd_sc_hd__nand2_1 _08822_ (.A(_03243_),
    .B(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__o21ba_1 _08823_ (.A1(_03179_),
    .A2(_03213_),
    .B1_N(_03212_),
    .X(_03246_));
 sky130_fd_sc_hd__nor2_1 _08824_ (.A(_03210_),
    .B(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__xnor2_1 _08825_ (.A(_03245_),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__o21ai_1 _08826_ (.A1(_01354_),
    .A2(_03248_),
    .B1(_01412_),
    .Y(_03249_));
 sky130_fd_sc_hd__a31o_1 _08827_ (.A1(_01355_),
    .A2(_03241_),
    .A3(_03242_),
    .B1(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__o211a_1 _08828_ (.A1(_02807_),
    .A2(_02845_),
    .B1(_02834_),
    .C1(_03250_),
    .X(_00383_));
 sky130_fd_sc_hd__nand2_1 _08829_ (.A(_03233_),
    .B(_03235_),
    .Y(_03251_));
 sky130_fd_sc_hd__a21o_1 _08830_ (.A1(_03229_),
    .A2(_03232_),
    .B1(_03228_),
    .X(_03252_));
 sky130_fd_sc_hd__xnor2_1 _08831_ (.A(_02817_),
    .B(\_225_[3] ),
    .Y(_03253_));
 sky130_fd_sc_hd__xnor2_2 _08832_ (.A(_02855_),
    .B(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__xnor2_1 _08833_ (.A(\_185_[13] ),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__xnor2_1 _08834_ (.A(_02064_),
    .B(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__nand2_1 _08835_ (.A(\_185_[12] ),
    .B(_03221_),
    .Y(_03257_));
 sky130_fd_sc_hd__o21a_1 _08836_ (.A1(_02071_),
    .A2(_03222_),
    .B1(_03257_),
    .X(_03258_));
 sky130_fd_sc_hd__xor2_1 _08837_ (.A(_03256_),
    .B(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__xnor2_1 _08838_ (.A(_02074_),
    .B(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__nor2_1 _08839_ (.A(_03223_),
    .B(_03225_),
    .Y(_03261_));
 sky130_fd_sc_hd__a21oi_1 _08840_ (.A1(_02048_),
    .A2(_03226_),
    .B1(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__xnor2_1 _08841_ (.A(_03260_),
    .B(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__a21o_1 _08842_ (.A1(\_228_[13] ),
    .A2(\_231_[13] ),
    .B1(_02811_),
    .X(_03264_));
 sky130_fd_sc_hd__o21a_1 _08843_ (.A1(\_228_[13] ),
    .A2(\_231_[13] ),
    .B1(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__xnor2_1 _08844_ (.A(_03263_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__xor2_1 _08845_ (.A(_03252_),
    .B(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__a21oi_1 _08846_ (.A1(_03251_),
    .A2(_03241_),
    .B1(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__a31o_1 _08847_ (.A1(_03251_),
    .A2(_03241_),
    .A3(_03267_),
    .B1(_01408_),
    .X(_03269_));
 sky130_fd_sc_hd__or2_1 _08848_ (.A(\_170_[13] ),
    .B(_02811_),
    .X(_03270_));
 sky130_fd_sc_hd__nand2_1 _08849_ (.A(\_170_[13] ),
    .B(_02811_),
    .Y(_03271_));
 sky130_fd_sc_hd__nand2_1 _08850_ (.A(_03270_),
    .B(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__o21ba_1 _08851_ (.A1(_03210_),
    .A2(_03246_),
    .B1_N(_03245_),
    .X(_03273_));
 sky130_fd_sc_hd__a21oi_1 _08852_ (.A1(\_170_[12] ),
    .A2(_02807_),
    .B1(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__xnor2_2 _08853_ (.A(_03272_),
    .B(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__nand2_1 _08854_ (.A(_02404_),
    .B(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__o211a_1 _08855_ (.A1(_03268_),
    .A2(_03269_),
    .B1(_03276_),
    .C1(_01439_),
    .X(_03277_));
 sky130_fd_sc_hd__a211o_1 _08856_ (.A1(_02811_),
    .A2(_03032_),
    .B1(_02861_),
    .C1(_03277_),
    .X(_00384_));
 sky130_fd_sc_hd__xnor2_1 _08857_ (.A(_02820_),
    .B(_02781_),
    .Y(_03278_));
 sky130_fd_sc_hd__xnor2_2 _08858_ (.A(_02858_),
    .B(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__xnor2_1 _08859_ (.A(\_185_[14] ),
    .B(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__xnor2_1 _08860_ (.A(_02124_),
    .B(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__nand2_1 _08861_ (.A(\_185_[13] ),
    .B(_03254_),
    .Y(_03282_));
 sky130_fd_sc_hd__o21a_1 _08862_ (.A1(_02064_),
    .A2(_03255_),
    .B1(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__xor2_1 _08863_ (.A(_03281_),
    .B(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__xnor2_1 _08864_ (.A(_02097_),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__nor2_1 _08865_ (.A(_03256_),
    .B(_03258_),
    .Y(_03286_));
 sky130_fd_sc_hd__a21oi_1 _08866_ (.A1(_02074_),
    .A2(_03259_),
    .B1(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__nor2_1 _08867_ (.A(_03285_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__and2_1 _08868_ (.A(_03285_),
    .B(_03287_),
    .X(_03289_));
 sky130_fd_sc_hd__or2_1 _08869_ (.A(_03288_),
    .B(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__a21o_1 _08870_ (.A1(\_228_[14] ),
    .A2(\_231_[14] ),
    .B1(_02814_),
    .X(_03291_));
 sky130_fd_sc_hd__o21a_1 _08871_ (.A1(\_228_[14] ),
    .A2(\_231_[14] ),
    .B1(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__xnor2_1 _08872_ (.A(_03290_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__or2b_1 _08873_ (.A(_03263_),
    .B_N(_03265_),
    .X(_03294_));
 sky130_fd_sc_hd__o21a_1 _08874_ (.A1(_03260_),
    .A2(_03262_),
    .B1(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__xor2_1 _08875_ (.A(_03293_),
    .B(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__nand2_1 _08876_ (.A(_03252_),
    .B(_03266_),
    .Y(_03297_));
 sky130_fd_sc_hd__nor2_1 _08877_ (.A(_03252_),
    .B(_03266_),
    .Y(_03298_));
 sky130_fd_sc_hd__a31o_1 _08878_ (.A1(_03251_),
    .A2(_03241_),
    .A3(_03297_),
    .B1(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__xor2_1 _08879_ (.A(_03296_),
    .B(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__nor2_1 _08880_ (.A(\_170_[14] ),
    .B(_02814_),
    .Y(_03301_));
 sky130_fd_sc_hd__nand2_1 _08881_ (.A(\_170_[14] ),
    .B(_02814_),
    .Y(_03302_));
 sky130_fd_sc_hd__and2b_1 _08882_ (.A_N(_03301_),
    .B(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__nand2_1 _08883_ (.A(_03244_),
    .B(_03271_),
    .Y(_03304_));
 sky130_fd_sc_hd__o21ai_2 _08884_ (.A1(_03273_),
    .A2(_03304_),
    .B1(_03270_),
    .Y(_03305_));
 sky130_fd_sc_hd__xor2_2 _08885_ (.A(_03303_),
    .B(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__nand2_1 _08886_ (.A(_02404_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__o211a_1 _08887_ (.A1(_02380_),
    .A2(_03300_),
    .B1(_03307_),
    .C1(_01439_),
    .X(_03308_));
 sky130_fd_sc_hd__a211o_1 _08888_ (.A1(_02814_),
    .A2(_03032_),
    .B1(_02861_),
    .C1(_03308_),
    .X(_00385_));
 sky130_fd_sc_hd__buf_6 _08889_ (.A(_01417_),
    .X(_03309_));
 sky130_fd_sc_hd__or2b_1 _08890_ (.A(_03295_),
    .B_N(_03293_),
    .X(_03310_));
 sky130_fd_sc_hd__or2_1 _08891_ (.A(_03296_),
    .B(_03299_),
    .X(_03311_));
 sky130_fd_sc_hd__and2b_1 _08892_ (.A_N(_03290_),
    .B(_03292_),
    .X(_03312_));
 sky130_fd_sc_hd__xnor2_1 _08893_ (.A(_02823_),
    .B(_02784_),
    .Y(_03313_));
 sky130_fd_sc_hd__xnor2_1 _08894_ (.A(_02862_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__xnor2_1 _08895_ (.A(\_185_[15] ),
    .B(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__xnor2_1 _08896_ (.A(_02117_),
    .B(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__nand2_1 _08897_ (.A(\_185_[14] ),
    .B(_03279_),
    .Y(_03317_));
 sky130_fd_sc_hd__o21a_1 _08898_ (.A1(_02124_),
    .A2(_03280_),
    .B1(_03317_),
    .X(_03318_));
 sky130_fd_sc_hd__xor2_1 _08899_ (.A(_03316_),
    .B(_03318_),
    .X(_03319_));
 sky130_fd_sc_hd__xnor2_1 _08900_ (.A(_02127_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__nor2_1 _08901_ (.A(_03281_),
    .B(_03283_),
    .Y(_03321_));
 sky130_fd_sc_hd__a21oi_1 _08902_ (.A1(_02097_),
    .A2(_03284_),
    .B1(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__nor2_1 _08903_ (.A(_03320_),
    .B(_03322_),
    .Y(_03323_));
 sky130_fd_sc_hd__nand2_1 _08904_ (.A(_03320_),
    .B(_03322_),
    .Y(_03324_));
 sky130_fd_sc_hd__or2b_1 _08905_ (.A(_03323_),
    .B_N(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__a21o_1 _08906_ (.A1(\_228_[15] ),
    .A2(\_231_[15] ),
    .B1(_02817_),
    .X(_03326_));
 sky130_fd_sc_hd__o21a_2 _08907_ (.A1(\_228_[15] ),
    .A2(\_231_[15] ),
    .B1(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__xnor2_1 _08908_ (.A(_03325_),
    .B(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__nor3_1 _08909_ (.A(_03288_),
    .B(_03312_),
    .C(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__o21a_1 _08910_ (.A1(_03288_),
    .A2(_03312_),
    .B1(_03328_),
    .X(_03330_));
 sky130_fd_sc_hd__nor2_1 _08911_ (.A(_03329_),
    .B(_03330_),
    .Y(_03331_));
 sky130_fd_sc_hd__and3_1 _08912_ (.A(_03310_),
    .B(_03311_),
    .C(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__a21oi_1 _08913_ (.A1(_03310_),
    .A2(_03311_),
    .B1(_03331_),
    .Y(_03333_));
 sky130_fd_sc_hd__nor2_1 _08914_ (.A(\_170_[15] ),
    .B(_02817_),
    .Y(_03334_));
 sky130_fd_sc_hd__and2_1 _08915_ (.A(\_170_[15] ),
    .B(_02817_),
    .X(_03335_));
 sky130_fd_sc_hd__nor2_1 _08916_ (.A(_03334_),
    .B(_03335_),
    .Y(_03336_));
 sky130_fd_sc_hd__o21ai_1 _08917_ (.A1(_03301_),
    .A2(_03305_),
    .B1(_03302_),
    .Y(_03337_));
 sky130_fd_sc_hd__xnor2_2 _08918_ (.A(_03336_),
    .B(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__nand2_1 _08919_ (.A(_01409_),
    .B(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__o311a_1 _08920_ (.A1(_01409_),
    .A2(_03332_),
    .A3(_03333_),
    .B1(_03339_),
    .C1(_01799_),
    .X(_03340_));
 sky130_fd_sc_hd__a211o_1 _08921_ (.A1(_02817_),
    .A2(_03032_),
    .B1(_03309_),
    .C1(_03340_),
    .X(_00386_));
 sky130_fd_sc_hd__nand2_1 _08922_ (.A(\_185_[15] ),
    .B(_03314_),
    .Y(_03341_));
 sky130_fd_sc_hd__or2_1 _08923_ (.A(_02117_),
    .B(_03315_),
    .X(_03342_));
 sky130_fd_sc_hd__xnor2_1 _08924_ (.A(_02827_),
    .B(_02787_),
    .Y(_03343_));
 sky130_fd_sc_hd__xnor2_1 _08925_ (.A(_02865_),
    .B(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__xnor2_1 _08926_ (.A(\_185_[16] ),
    .B(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__xnor2_1 _08927_ (.A(_02151_),
    .B(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__a21o_1 _08928_ (.A1(_03341_),
    .A2(_03342_),
    .B1(_03346_),
    .X(_03347_));
 sky130_fd_sc_hd__nand3_1 _08929_ (.A(_03341_),
    .B(_03342_),
    .C(_03346_),
    .Y(_03348_));
 sky130_fd_sc_hd__and3_1 _08930_ (.A(_02161_),
    .B(_03347_),
    .C(_03348_),
    .X(_03349_));
 sky130_fd_sc_hd__a21oi_1 _08931_ (.A1(_03347_),
    .A2(_03348_),
    .B1(_02161_),
    .Y(_03350_));
 sky130_fd_sc_hd__or2_1 _08932_ (.A(_03349_),
    .B(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__nor2_1 _08933_ (.A(_03316_),
    .B(_03318_),
    .Y(_03352_));
 sky130_fd_sc_hd__a21oi_2 _08934_ (.A1(_02127_),
    .A2(_03319_),
    .B1(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__xnor2_1 _08935_ (.A(_03351_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__a21o_1 _08936_ (.A1(\_228_[16] ),
    .A2(\_231_[16] ),
    .B1(_02820_),
    .X(_03355_));
 sky130_fd_sc_hd__o21a_1 _08937_ (.A1(\_228_[16] ),
    .A2(\_231_[16] ),
    .B1(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__xnor2_1 _08938_ (.A(_03354_),
    .B(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__a21oi_2 _08939_ (.A1(_03324_),
    .A2(_03327_),
    .B1(_03323_),
    .Y(_03358_));
 sky130_fd_sc_hd__xnor2_2 _08940_ (.A(_03357_),
    .B(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__or3_1 _08941_ (.A(_03296_),
    .B(_03329_),
    .C(_03330_),
    .X(_03360_));
 sky130_fd_sc_hd__a21o_1 _08942_ (.A1(_03251_),
    .A2(_03297_),
    .B1(_03298_),
    .X(_03361_));
 sky130_fd_sc_hd__inv_2 _08943_ (.A(_03330_),
    .Y(_03362_));
 sky130_fd_sc_hd__o221a_1 _08944_ (.A1(_03310_),
    .A2(_03329_),
    .B1(_03360_),
    .B2(_03361_),
    .C1(_03362_),
    .X(_03363_));
 sky130_fd_sc_hd__nand2_1 _08945_ (.A(_03236_),
    .B(_03267_),
    .Y(_03364_));
 sky130_fd_sc_hd__or3_1 _08946_ (.A(_03239_),
    .B(_03364_),
    .C(_03360_),
    .X(_03365_));
 sky130_fd_sc_hd__a2111o_1 _08947_ (.A1(_03095_),
    .A2(_03099_),
    .B1(_03238_),
    .C1(_03364_),
    .D1(_03360_),
    .X(_03366_));
 sky130_fd_sc_hd__and3_1 _08948_ (.A(_03363_),
    .B(_03365_),
    .C(_03366_),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_2 _08949_ (.A(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__xnor2_1 _08950_ (.A(_03359_),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__or2_1 _08951_ (.A(\_170_[16] ),
    .B(_02820_),
    .X(_03370_));
 sky130_fd_sc_hd__nand2_1 _08952_ (.A(\_170_[16] ),
    .B(_02820_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand2_2 _08953_ (.A(_03370_),
    .B(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__o211a_1 _08954_ (.A1(\_170_[15] ),
    .A2(_02817_),
    .B1(_02814_),
    .C1(\_170_[14] ),
    .X(_03373_));
 sky130_fd_sc_hd__o2111a_1 _08955_ (.A1(_03273_),
    .A2(_03304_),
    .B1(_03336_),
    .C1(_03270_),
    .D1(_03303_),
    .X(_03374_));
 sky130_fd_sc_hd__nor3_4 _08956_ (.A(_03335_),
    .B(_03373_),
    .C(_03374_),
    .Y(_03375_));
 sky130_fd_sc_hd__xnor2_2 _08957_ (.A(_03372_),
    .B(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__nand2_1 _08958_ (.A(_02404_),
    .B(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__o211a_1 _08959_ (.A1(_02380_),
    .A2(_03369_),
    .B1(_03377_),
    .C1(_01439_),
    .X(_03378_));
 sky130_fd_sc_hd__a211o_1 _08960_ (.A1(_02820_),
    .A2(_03032_),
    .B1(_03309_),
    .C1(_03378_),
    .X(_00387_));
 sky130_fd_sc_hd__buf_6 _08961_ (.A(_02833_),
    .X(_03379_));
 sky130_fd_sc_hd__nor2_1 _08962_ (.A(_03351_),
    .B(_03353_),
    .Y(_03380_));
 sky130_fd_sc_hd__and2b_1 _08963_ (.A_N(_03354_),
    .B(_03356_),
    .X(_03381_));
 sky130_fd_sc_hd__xnor2_1 _08964_ (.A(_02830_),
    .B(_02790_),
    .Y(_03382_));
 sky130_fd_sc_hd__xnor2_1 _08965_ (.A(_02868_),
    .B(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__xnor2_1 _08966_ (.A(\_185_[17] ),
    .B(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__xnor2_1 _08967_ (.A(_02205_),
    .B(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__nand2_1 _08968_ (.A(\_185_[16] ),
    .B(_03344_),
    .Y(_03386_));
 sky130_fd_sc_hd__o21a_1 _08969_ (.A1(_02151_),
    .A2(_03345_),
    .B1(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__xor2_1 _08970_ (.A(_03385_),
    .B(_03387_),
    .X(_03388_));
 sky130_fd_sc_hd__xnor2_1 _08971_ (.A(_02192_),
    .B(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__a21boi_2 _08972_ (.A1(_02161_),
    .A2(_03348_),
    .B1_N(_03347_),
    .Y(_03390_));
 sky130_fd_sc_hd__xnor2_1 _08973_ (.A(_03389_),
    .B(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__a21o_1 _08974_ (.A1(\_228_[17] ),
    .A2(\_231_[17] ),
    .B1(_02823_),
    .X(_03392_));
 sky130_fd_sc_hd__o21a_1 _08975_ (.A1(\_228_[17] ),
    .A2(\_231_[17] ),
    .B1(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__xnor2_1 _08976_ (.A(_03391_),
    .B(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__o21ai_1 _08977_ (.A1(_03380_),
    .A2(_03381_),
    .B1(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__nor3_1 _08978_ (.A(_03380_),
    .B(_03381_),
    .C(_03394_),
    .Y(_03396_));
 sky130_fd_sc_hd__inv_2 _08979_ (.A(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_1 _08980_ (.A(_03395_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__inv_2 _08981_ (.A(_03359_),
    .Y(_03399_));
 sky130_fd_sc_hd__or2b_1 _08982_ (.A(_03358_),
    .B_N(_03357_),
    .X(_03400_));
 sky130_fd_sc_hd__o21ai_1 _08983_ (.A1(_03399_),
    .A2(_03368_),
    .B1(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__xnor2_1 _08984_ (.A(_03398_),
    .B(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__nand2_1 _08985_ (.A(\_170_[17] ),
    .B(_02823_),
    .Y(_03403_));
 sky130_fd_sc_hd__or2_1 _08986_ (.A(\_170_[17] ),
    .B(_02823_),
    .X(_03404_));
 sky130_fd_sc_hd__nand2_1 _08987_ (.A(_03403_),
    .B(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__o21ai_2 _08988_ (.A1(_03372_),
    .A2(_03375_),
    .B1(_03371_),
    .Y(_03406_));
 sky130_fd_sc_hd__xor2_2 _08989_ (.A(_03405_),
    .B(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__nor2_1 _08990_ (.A(_01778_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__a211o_1 _08991_ (.A1(_01520_),
    .A2(_03402_),
    .B1(_03408_),
    .C1(_02355_),
    .X(_03409_));
 sky130_fd_sc_hd__o211a_1 _08992_ (.A1(_02823_),
    .A2(_02845_),
    .B1(_03379_),
    .C1(_03409_),
    .X(_00388_));
 sky130_fd_sc_hd__nor2_1 _08993_ (.A(_03389_),
    .B(_03390_),
    .Y(_03410_));
 sky130_fd_sc_hd__and2b_1 _08994_ (.A_N(_03391_),
    .B(_03393_),
    .X(_03411_));
 sky130_fd_sc_hd__xnor2_1 _08995_ (.A(_02835_),
    .B(_02794_),
    .Y(_03412_));
 sky130_fd_sc_hd__xnor2_2 _08996_ (.A(_02871_),
    .B(_03412_),
    .Y(_03413_));
 sky130_fd_sc_hd__xnor2_1 _08997_ (.A(\_185_[18] ),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__xnor2_1 _08998_ (.A(_02249_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand2_1 _08999_ (.A(\_185_[17] ),
    .B(_03383_),
    .Y(_03416_));
 sky130_fd_sc_hd__o21a_1 _09000_ (.A1(_02205_),
    .A2(_03384_),
    .B1(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__xor2_1 _09001_ (.A(_03415_),
    .B(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__xnor2_1 _09002_ (.A(_02216_),
    .B(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__nor2_1 _09003_ (.A(_03385_),
    .B(_03387_),
    .Y(_03420_));
 sky130_fd_sc_hd__a21oi_1 _09004_ (.A1(_02192_),
    .A2(_03388_),
    .B1(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hd__xnor2_1 _09005_ (.A(_03419_),
    .B(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__a21o_1 _09006_ (.A1(\_228_[18] ),
    .A2(\_231_[18] ),
    .B1(_02827_),
    .X(_03423_));
 sky130_fd_sc_hd__o21a_1 _09007_ (.A1(\_228_[18] ),
    .A2(\_231_[18] ),
    .B1(_03423_),
    .X(_03424_));
 sky130_fd_sc_hd__xnor2_1 _09008_ (.A(_03422_),
    .B(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__o21ai_1 _09009_ (.A1(_03410_),
    .A2(_03411_),
    .B1(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__or3_1 _09010_ (.A(_03410_),
    .B(_03411_),
    .C(_03425_),
    .X(_03427_));
 sky130_fd_sc_hd__and2_1 _09011_ (.A(_03426_),
    .B(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__nand3b_1 _09012_ (.A_N(_03396_),
    .B(_03359_),
    .C(_03395_),
    .Y(_03429_));
 sky130_fd_sc_hd__a21oi_1 _09013_ (.A1(_03400_),
    .A2(_03395_),
    .B1(_03396_),
    .Y(_03430_));
 sky130_fd_sc_hd__o21bai_1 _09014_ (.A1(_03368_),
    .A2(_03429_),
    .B1_N(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_1 _09015_ (.A(_03428_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__o21a_1 _09016_ (.A1(_03428_),
    .A2(_03431_),
    .B1(_01523_),
    .X(_03433_));
 sky130_fd_sc_hd__nor2_1 _09017_ (.A(\_170_[18] ),
    .B(_02827_),
    .Y(_03434_));
 sky130_fd_sc_hd__and2_1 _09018_ (.A(\_170_[18] ),
    .B(_02827_),
    .X(_03435_));
 sky130_fd_sc_hd__nor2_1 _09019_ (.A(_03434_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__a21bo_1 _09020_ (.A1(_03404_),
    .A2(_03406_),
    .B1_N(_03403_),
    .X(_03437_));
 sky130_fd_sc_hd__xnor2_1 _09021_ (.A(_03436_),
    .B(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__nor2_1 _09022_ (.A(_01778_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__a211o_1 _09023_ (.A1(_03432_),
    .A2(_03433_),
    .B1(_03439_),
    .C1(_02355_),
    .X(_03440_));
 sky130_fd_sc_hd__o211a_1 _09024_ (.A1(_02827_),
    .A2(_01426_),
    .B1(_03379_),
    .C1(_03440_),
    .X(_00389_));
 sky130_fd_sc_hd__nor2_1 _09025_ (.A(_03419_),
    .B(_03421_),
    .Y(_03441_));
 sky130_fd_sc_hd__and2b_1 _09026_ (.A_N(_03422_),
    .B(_03424_),
    .X(_03442_));
 sky130_fd_sc_hd__xnor2_1 _09027_ (.A(_02797_),
    .B(_02768_),
    .Y(_03443_));
 sky130_fd_sc_hd__xnor2_2 _09028_ (.A(_02839_),
    .B(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__xnor2_1 _09029_ (.A(\_185_[19] ),
    .B(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__xnor2_1 _09030_ (.A(_02242_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_1 _09031_ (.A(\_185_[18] ),
    .B(_03413_),
    .Y(_03447_));
 sky130_fd_sc_hd__o21ai_1 _09032_ (.A1(_02249_),
    .A2(_03414_),
    .B1(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hd__xnor2_1 _09033_ (.A(_03446_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__xnor2_1 _09034_ (.A(_02252_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__nor2_1 _09035_ (.A(_03415_),
    .B(_03417_),
    .Y(_03451_));
 sky130_fd_sc_hd__a21oi_1 _09036_ (.A1(_02216_),
    .A2(_03418_),
    .B1(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__xnor2_1 _09037_ (.A(_03450_),
    .B(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__a21o_1 _09038_ (.A1(\_228_[19] ),
    .A2(\_231_[19] ),
    .B1(_02830_),
    .X(_03454_));
 sky130_fd_sc_hd__o21a_1 _09039_ (.A1(\_228_[19] ),
    .A2(\_231_[19] ),
    .B1(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__xnor2_1 _09040_ (.A(_03453_),
    .B(_03455_),
    .Y(_03456_));
 sky130_fd_sc_hd__nor3_1 _09041_ (.A(_03441_),
    .B(_03442_),
    .C(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__o21ai_1 _09042_ (.A1(_03441_),
    .A2(_03442_),
    .B1(_03456_),
    .Y(_03458_));
 sky130_fd_sc_hd__and2b_1 _09043_ (.A_N(_03457_),
    .B(_03458_),
    .X(_03459_));
 sky130_fd_sc_hd__and3_1 _09044_ (.A(_03426_),
    .B(_03432_),
    .C(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__a21oi_1 _09045_ (.A1(_03426_),
    .A2(_03432_),
    .B1(_03459_),
    .Y(_03461_));
 sky130_fd_sc_hd__xor2_2 _09046_ (.A(\_170_[19] ),
    .B(_02830_),
    .X(_03462_));
 sky130_fd_sc_hd__a21oi_1 _09047_ (.A1(_03436_),
    .A2(_03437_),
    .B1(_03435_),
    .Y(_03463_));
 sky130_fd_sc_hd__xor2_2 _09048_ (.A(_03462_),
    .B(_03463_),
    .X(_03464_));
 sky130_fd_sc_hd__nand2_1 _09049_ (.A(_01409_),
    .B(_03464_),
    .Y(_03465_));
 sky130_fd_sc_hd__o311a_1 _09050_ (.A1(_01409_),
    .A2(_03460_),
    .A3(_03461_),
    .B1(_03465_),
    .C1(_01799_),
    .X(_03466_));
 sky130_fd_sc_hd__a211o_1 _09051_ (.A1(_02830_),
    .A2(_03032_),
    .B1(_03309_),
    .C1(_03466_),
    .X(_00390_));
 sky130_fd_sc_hd__nor2_1 _09052_ (.A(\_170_[20] ),
    .B(_02835_),
    .Y(_03467_));
 sky130_fd_sc_hd__nand2_1 _09053_ (.A(\_170_[20] ),
    .B(_02835_),
    .Y(_03468_));
 sky130_fd_sc_hd__or2b_1 _09054_ (.A(_03467_),
    .B_N(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__or4bb_1 _09055_ (.A(_03372_),
    .B(_03405_),
    .C_N(_03436_),
    .D_N(_03462_),
    .X(_03470_));
 sky130_fd_sc_hd__nand2_1 _09056_ (.A(_03371_),
    .B(_03403_),
    .Y(_03471_));
 sky130_fd_sc_hd__and4_1 _09057_ (.A(_03404_),
    .B(_03436_),
    .C(_03471_),
    .D(_03462_),
    .X(_03472_));
 sky130_fd_sc_hd__o21a_1 _09058_ (.A1(\_170_[19] ),
    .A2(_02830_),
    .B1(_03435_),
    .X(_03473_));
 sky130_fd_sc_hd__a211oi_1 _09059_ (.A1(\_170_[19] ),
    .A2(_02830_),
    .B1(_03472_),
    .C1(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__o21ai_1 _09060_ (.A1(_03375_),
    .A2(_03470_),
    .B1(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__and2b_1 _09061_ (.A_N(_03469_),
    .B(_03475_),
    .X(_03476_));
 sky130_fd_sc_hd__and2b_1 _09062_ (.A_N(_03475_),
    .B(_03469_),
    .X(_03477_));
 sky130_fd_sc_hd__nor2_1 _09063_ (.A(_03476_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__nor2_1 _09064_ (.A(_03450_),
    .B(_03452_),
    .Y(_03479_));
 sky130_fd_sc_hd__and2b_1 _09065_ (.A_N(_03453_),
    .B(_03455_),
    .X(_03480_));
 sky130_fd_sc_hd__or2b_1 _09066_ (.A(_03446_),
    .B_N(_03448_),
    .X(_03481_));
 sky130_fd_sc_hd__nand2_1 _09067_ (.A(_02252_),
    .B(_03449_),
    .Y(_03482_));
 sky130_fd_sc_hd__xnor2_1 _09068_ (.A(_02801_),
    .B(_02772_),
    .Y(_03483_));
 sky130_fd_sc_hd__xnor2_2 _09069_ (.A(_02842_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__xor2_1 _09070_ (.A(\_185_[20] ),
    .B(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__xnor2_1 _09071_ (.A(_02262_),
    .B(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__nand2_1 _09072_ (.A(\_185_[19] ),
    .B(_03444_),
    .Y(_03487_));
 sky130_fd_sc_hd__o21ai_1 _09073_ (.A1(_02242_),
    .A2(_03445_),
    .B1(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__xnor2_1 _09074_ (.A(_03486_),
    .B(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__xnor2_1 _09075_ (.A(_02271_),
    .B(_03489_),
    .Y(_03490_));
 sky130_fd_sc_hd__a21oi_1 _09076_ (.A1(_03481_),
    .A2(_03482_),
    .B1(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__and3_1 _09077_ (.A(_03481_),
    .B(_03482_),
    .C(_03490_),
    .X(_03492_));
 sky130_fd_sc_hd__or2_1 _09078_ (.A(_03491_),
    .B(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__a21o_1 _09079_ (.A1(\_228_[20] ),
    .A2(\_231_[20] ),
    .B1(_02835_),
    .X(_03494_));
 sky130_fd_sc_hd__o21a_1 _09080_ (.A1(\_228_[20] ),
    .A2(\_231_[20] ),
    .B1(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__xnor2_1 _09081_ (.A(_03493_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__o21ai_1 _09082_ (.A1(_03479_),
    .A2(_03480_),
    .B1(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__or3_1 _09083_ (.A(_03479_),
    .B(_03480_),
    .C(_03496_),
    .X(_03498_));
 sky130_fd_sc_hd__and2_1 _09084_ (.A(_03497_),
    .B(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__nand2_1 _09085_ (.A(_03428_),
    .B(_03459_),
    .Y(_03500_));
 sky130_fd_sc_hd__or2_1 _09086_ (.A(_03429_),
    .B(_03500_),
    .X(_03501_));
 sky130_fd_sc_hd__or2b_1 _09087_ (.A(_03500_),
    .B_N(_03430_),
    .X(_03502_));
 sky130_fd_sc_hd__o211a_1 _09088_ (.A1(_03426_),
    .A2(_03457_),
    .B1(_03458_),
    .C1(_03502_),
    .X(_03503_));
 sky130_fd_sc_hd__o21ai_2 _09089_ (.A1(_03368_),
    .A2(_03501_),
    .B1(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__o21ai_1 _09090_ (.A1(_03499_),
    .A2(_03504_),
    .B1(_01523_),
    .Y(_03505_));
 sky130_fd_sc_hd__a21oi_1 _09091_ (.A1(_03499_),
    .A2(_03504_),
    .B1(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__a211o_1 _09092_ (.A1(_01856_),
    .A2(_03478_),
    .B1(_03506_),
    .C1(_01495_),
    .X(_03507_));
 sky130_fd_sc_hd__o211a_1 _09093_ (.A1(_02835_),
    .A2(_01426_),
    .B1(_03379_),
    .C1(_03507_),
    .X(_00391_));
 sky130_fd_sc_hd__nand2_1 _09094_ (.A(\_170_[21] ),
    .B(_02839_),
    .Y(_03508_));
 sky130_fd_sc_hd__or2_1 _09095_ (.A(\_170_[21] ),
    .B(_02839_),
    .X(_03509_));
 sky130_fd_sc_hd__nand2_1 _09096_ (.A(_03508_),
    .B(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__a21o_1 _09097_ (.A1(\_170_[20] ),
    .A2(_02835_),
    .B1(_03476_),
    .X(_03511_));
 sky130_fd_sc_hd__xnor2_2 _09098_ (.A(_03510_),
    .B(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__and2b_1 _09099_ (.A_N(_03493_),
    .B(_03495_),
    .X(_03513_));
 sky130_fd_sc_hd__or2b_1 _09100_ (.A(_03486_),
    .B_N(_03488_),
    .X(_03514_));
 sky130_fd_sc_hd__nand2_1 _09101_ (.A(_02271_),
    .B(_03489_),
    .Y(_03515_));
 sky130_fd_sc_hd__nand2_1 _09102_ (.A(_03514_),
    .B(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__or2_1 _09103_ (.A(\_185_[20] ),
    .B(_03484_),
    .X(_03517_));
 sky130_fd_sc_hd__and2_1 _09104_ (.A(\_185_[20] ),
    .B(_03484_),
    .X(_03518_));
 sky130_fd_sc_hd__a21oi_1 _09105_ (.A1(_02262_),
    .A2(_03517_),
    .B1(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__xnor2_1 _09106_ (.A(_02804_),
    .B(_02776_),
    .Y(_03520_));
 sky130_fd_sc_hd__xnor2_1 _09107_ (.A(_02846_),
    .B(_03520_),
    .Y(_03521_));
 sky130_fd_sc_hd__nand2_1 _09108_ (.A(\_185_[21] ),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__or2_1 _09109_ (.A(\_185_[21] ),
    .B(_03521_),
    .X(_03523_));
 sky130_fd_sc_hd__nand2_1 _09110_ (.A(_03522_),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__xnor2_1 _09111_ (.A(_02323_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__xor2_1 _09112_ (.A(_03519_),
    .B(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__xnor2_1 _09113_ (.A(_02311_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__xnor2_1 _09114_ (.A(_03516_),
    .B(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__a21o_1 _09115_ (.A1(\_228_[21] ),
    .A2(\_231_[21] ),
    .B1(_02839_),
    .X(_03529_));
 sky130_fd_sc_hd__o21a_1 _09116_ (.A1(\_228_[21] ),
    .A2(\_231_[21] ),
    .B1(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__xor2_1 _09117_ (.A(_03528_),
    .B(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__o21ai_1 _09118_ (.A1(_03491_),
    .A2(_03513_),
    .B1(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__or3_1 _09119_ (.A(_03491_),
    .B(_03513_),
    .C(_03531_),
    .X(_03533_));
 sky130_fd_sc_hd__and2_1 _09120_ (.A(_03532_),
    .B(_03533_),
    .X(_03534_));
 sky130_fd_sc_hd__a21bo_1 _09121_ (.A1(_03499_),
    .A2(_03504_),
    .B1_N(_03497_),
    .X(_03535_));
 sky130_fd_sc_hd__nand2_1 _09122_ (.A(_03534_),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__o211a_1 _09123_ (.A1(_03534_),
    .A2(_03535_),
    .B1(_03536_),
    .C1(_01523_),
    .X(_03537_));
 sky130_fd_sc_hd__a211o_1 _09124_ (.A1(_01428_),
    .A2(_03512_),
    .B1(_03537_),
    .C1(_01495_),
    .X(_03538_));
 sky130_fd_sc_hd__o211a_1 _09125_ (.A1(_02839_),
    .A2(_01426_),
    .B1(_03379_),
    .C1(_03538_),
    .X(_00392_));
 sky130_fd_sc_hd__nor2_1 _09126_ (.A(\_170_[22] ),
    .B(_02842_),
    .Y(_03539_));
 sky130_fd_sc_hd__and2_1 _09127_ (.A(\_170_[22] ),
    .B(_02842_),
    .X(_03540_));
 sky130_fd_sc_hd__nor2_1 _09128_ (.A(_03539_),
    .B(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__nand2_1 _09129_ (.A(_03468_),
    .B(_03508_),
    .Y(_03542_));
 sky130_fd_sc_hd__o21a_1 _09130_ (.A1(_03476_),
    .A2(_03542_),
    .B1(_03509_),
    .X(_03543_));
 sky130_fd_sc_hd__xnor2_2 _09131_ (.A(_03541_),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__a21oi_1 _09132_ (.A1(_03514_),
    .A2(_03515_),
    .B1(_03527_),
    .Y(_03545_));
 sky130_fd_sc_hd__and2_1 _09133_ (.A(_03528_),
    .B(_03530_),
    .X(_03546_));
 sky130_fd_sc_hd__xnor2_1 _09134_ (.A(_02807_),
    .B(\_225_[3] ),
    .Y(_03547_));
 sky130_fd_sc_hd__xnor2_2 _09135_ (.A(_02849_),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__xnor2_1 _09136_ (.A(\_185_[22] ),
    .B(_03548_),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_1 _09137_ (.A(_02327_),
    .B(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__or2_1 _09138_ (.A(_02327_),
    .B(_03549_),
    .X(_03551_));
 sky130_fd_sc_hd__nand2_1 _09139_ (.A(_03550_),
    .B(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__o21ai_1 _09140_ (.A1(_02323_),
    .A2(_03524_),
    .B1(_03522_),
    .Y(_03553_));
 sky130_fd_sc_hd__xnor2_1 _09141_ (.A(_03552_),
    .B(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__xnor2_1 _09142_ (.A(_02337_),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__nor2_1 _09143_ (.A(_03519_),
    .B(_03525_),
    .Y(_03556_));
 sky130_fd_sc_hd__a21o_1 _09144_ (.A1(_02311_),
    .A2(_03526_),
    .B1(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__xor2_1 _09145_ (.A(_03555_),
    .B(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__a21o_1 _09146_ (.A1(\_228_[22] ),
    .A2(\_231_[22] ),
    .B1(_02842_),
    .X(_03559_));
 sky130_fd_sc_hd__o21a_1 _09147_ (.A1(\_228_[22] ),
    .A2(\_231_[22] ),
    .B1(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__xnor2_1 _09148_ (.A(_03558_),
    .B(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__o21ai_1 _09149_ (.A1(_03545_),
    .A2(_03546_),
    .B1(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__or3_1 _09150_ (.A(_03545_),
    .B(_03546_),
    .C(_03561_),
    .X(_03563_));
 sky130_fd_sc_hd__and2_1 _09151_ (.A(_03562_),
    .B(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__a21bo_1 _09152_ (.A1(_03497_),
    .A2(_03532_),
    .B1_N(_03533_),
    .X(_03565_));
 sky130_fd_sc_hd__inv_2 _09153_ (.A(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__a31o_1 _09154_ (.A1(_03499_),
    .A2(_03504_),
    .A3(_03534_),
    .B1(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__xnor2_1 _09155_ (.A(_03564_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__mux2_1 _09156_ (.A0(_03544_),
    .A1(_03568_),
    .S(_01354_),
    .X(_03569_));
 sky130_fd_sc_hd__nand2_1 _09157_ (.A(_01421_),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__o211a_1 _09158_ (.A1(_02842_),
    .A2(_01426_),
    .B1(_03379_),
    .C1(_03570_),
    .X(_00393_));
 sky130_fd_sc_hd__and2b_1 _09159_ (.A_N(_03555_),
    .B(_03557_),
    .X(_03571_));
 sky130_fd_sc_hd__and2b_1 _09160_ (.A_N(_03558_),
    .B(_03560_),
    .X(_03572_));
 sky130_fd_sc_hd__nand2_1 _09161_ (.A(\_185_[22] ),
    .B(_03548_),
    .Y(_03573_));
 sky130_fd_sc_hd__xnor2_1 _09162_ (.A(_02811_),
    .B(_02781_),
    .Y(_03574_));
 sky130_fd_sc_hd__xnor2_1 _09163_ (.A(_02852_),
    .B(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__xnor2_1 _09164_ (.A(\_185_[23] ),
    .B(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__xor2_1 _09165_ (.A(_02362_),
    .B(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__a21o_1 _09166_ (.A1(_03573_),
    .A2(_03551_),
    .B1(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__nand3_1 _09167_ (.A(_03573_),
    .B(_03551_),
    .C(_03577_),
    .Y(_03579_));
 sky130_fd_sc_hd__and2_1 _09168_ (.A(_03578_),
    .B(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__xnor2_1 _09169_ (.A(_02371_),
    .B(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__a32o_1 _09170_ (.A1(_03550_),
    .A2(_03551_),
    .A3(_03553_),
    .B1(_03554_),
    .B2(_02337_),
    .X(_03582_));
 sky130_fd_sc_hd__xor2_1 _09171_ (.A(_03581_),
    .B(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__a21o_1 _09172_ (.A1(\_228_[23] ),
    .A2(\_231_[23] ),
    .B1(_02846_),
    .X(_03584_));
 sky130_fd_sc_hd__o21ai_2 _09173_ (.A1(\_228_[23] ),
    .A2(\_231_[23] ),
    .B1(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__xor2_1 _09174_ (.A(_03583_),
    .B(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__nor3_1 _09175_ (.A(_03571_),
    .B(_03572_),
    .C(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__o21ai_1 _09176_ (.A1(_03571_),
    .A2(_03572_),
    .B1(_03586_),
    .Y(_03588_));
 sky130_fd_sc_hd__and2b_1 _09177_ (.A_N(_03587_),
    .B(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__a21bo_1 _09178_ (.A1(_03564_),
    .A2(_03567_),
    .B1_N(_03562_),
    .X(_03590_));
 sky130_fd_sc_hd__nand2_1 _09179_ (.A(_03589_),
    .B(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__o21a_1 _09180_ (.A1(_03589_),
    .A2(_03590_),
    .B1(_01354_),
    .X(_03592_));
 sky130_fd_sc_hd__xor2_2 _09181_ (.A(\_170_[23] ),
    .B(_02846_),
    .X(_03593_));
 sky130_fd_sc_hd__a21o_1 _09182_ (.A1(_03541_),
    .A2(_03543_),
    .B1(_03540_),
    .X(_03594_));
 sky130_fd_sc_hd__xor2_2 _09183_ (.A(_03593_),
    .B(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__a21o_1 _09184_ (.A1(_01923_),
    .A2(_03595_),
    .B1(_02002_),
    .X(_03596_));
 sky130_fd_sc_hd__a21o_1 _09185_ (.A1(_03591_),
    .A2(_03592_),
    .B1(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__o211a_1 _09186_ (.A1(_02846_),
    .A2(_01426_),
    .B1(_03379_),
    .C1(_03597_),
    .X(_00394_));
 sky130_fd_sc_hd__or2_1 _09187_ (.A(\_170_[24] ),
    .B(_02849_),
    .X(_03598_));
 sky130_fd_sc_hd__nand2_1 _09188_ (.A(\_170_[24] ),
    .B(_02849_),
    .Y(_03599_));
 sky130_fd_sc_hd__nand2_1 _09189_ (.A(_03598_),
    .B(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__or4bb_1 _09190_ (.A(_03469_),
    .B(_03510_),
    .C_N(_03541_),
    .D_N(_03593_),
    .X(_03601_));
 sky130_fd_sc_hd__o21bai_1 _09191_ (.A1(_03467_),
    .A2(_03474_),
    .B1_N(_03542_),
    .Y(_03602_));
 sky130_fd_sc_hd__a21o_1 _09192_ (.A1(_03509_),
    .A2(_03602_),
    .B1(_03540_),
    .X(_03603_));
 sky130_fd_sc_hd__o221a_1 _09193_ (.A1(\_170_[23] ),
    .A2(_02846_),
    .B1(_02842_),
    .B2(\_170_[22] ),
    .C1(_03603_),
    .X(_03604_));
 sky130_fd_sc_hd__a21oi_1 _09194_ (.A1(\_170_[23] ),
    .A2(_02846_),
    .B1(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__o31a_1 _09195_ (.A1(_03375_),
    .A2(_03470_),
    .A3(_03601_),
    .B1(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__xor2_2 _09196_ (.A(_03600_),
    .B(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__nand2_1 _09197_ (.A(\_185_[23] ),
    .B(_03575_),
    .Y(_03608_));
 sky130_fd_sc_hd__inv_2 _09198_ (.A(_03576_),
    .Y(_03609_));
 sky130_fd_sc_hd__nand2_1 _09199_ (.A(_02362_),
    .B(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__xnor2_1 _09200_ (.A(_02814_),
    .B(_02784_),
    .Y(_03611_));
 sky130_fd_sc_hd__xnor2_1 _09201_ (.A(_02855_),
    .B(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__xnor2_1 _09202_ (.A(\_185_[24] ),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__xor2_1 _09203_ (.A(_02383_),
    .B(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__a21o_1 _09204_ (.A1(_03608_),
    .A2(_03610_),
    .B1(_03614_),
    .X(_03615_));
 sky130_fd_sc_hd__nand3_1 _09205_ (.A(_03608_),
    .B(_03610_),
    .C(_03614_),
    .Y(_03616_));
 sky130_fd_sc_hd__and2_1 _09206_ (.A(_03615_),
    .B(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__or2_1 _09207_ (.A(_02392_),
    .B(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__nand2_1 _09208_ (.A(_02392_),
    .B(_03617_),
    .Y(_03619_));
 sky130_fd_sc_hd__nand2_1 _09209_ (.A(_03618_),
    .B(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__a21bo_1 _09210_ (.A1(_02371_),
    .A2(_03580_),
    .B1_N(_03578_),
    .X(_03621_));
 sky130_fd_sc_hd__xor2_1 _09211_ (.A(_03620_),
    .B(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__a21o_1 _09212_ (.A1(\_228_[24] ),
    .A2(\_231_[24] ),
    .B1(_02849_),
    .X(_03623_));
 sky130_fd_sc_hd__o21a_1 _09213_ (.A1(\_228_[24] ),
    .A2(\_231_[24] ),
    .B1(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__xnor2_1 _09214_ (.A(_03622_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__and2b_1 _09215_ (.A_N(_03581_),
    .B(_03582_),
    .X(_03626_));
 sky130_fd_sc_hd__o21ba_1 _09216_ (.A1(_03583_),
    .A2(_03585_),
    .B1_N(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__xnor2_1 _09217_ (.A(_03625_),
    .B(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__nand2_1 _09218_ (.A(_03564_),
    .B(_03589_),
    .Y(_03629_));
 sky130_fd_sc_hd__o221a_1 _09219_ (.A1(_03562_),
    .A2(_03587_),
    .B1(_03629_),
    .B2(_03565_),
    .C1(_03588_),
    .X(_03630_));
 sky130_fd_sc_hd__nand2_1 _09220_ (.A(_03499_),
    .B(_03534_),
    .Y(_03631_));
 sky130_fd_sc_hd__or3_1 _09221_ (.A(_03501_),
    .B(_03631_),
    .C(_03629_),
    .X(_03632_));
 sky130_fd_sc_hd__o32a_1 _09222_ (.A1(_03503_),
    .A2(_03631_),
    .A3(_03629_),
    .B1(_03632_),
    .B2(_03368_),
    .X(_03633_));
 sky130_fd_sc_hd__nand2_1 _09223_ (.A(_03630_),
    .B(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hd__nand2_1 _09224_ (.A(_03628_),
    .B(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__o211a_1 _09225_ (.A1(_03628_),
    .A2(_03634_),
    .B1(_03635_),
    .C1(_01523_),
    .X(_03636_));
 sky130_fd_sc_hd__a211o_1 _09226_ (.A1(_01428_),
    .A2(_03607_),
    .B1(_03636_),
    .C1(_01495_),
    .X(_03637_));
 sky130_fd_sc_hd__o211a_1 _09227_ (.A1(_02849_),
    .A2(_01426_),
    .B1(_03379_),
    .C1(_03637_),
    .X(_00395_));
 sky130_fd_sc_hd__and2b_1 _09228_ (.A_N(_03620_),
    .B(_03621_),
    .X(_03638_));
 sky130_fd_sc_hd__and2b_1 _09229_ (.A_N(_03622_),
    .B(_03624_),
    .X(_03639_));
 sky130_fd_sc_hd__nand2_1 _09230_ (.A(\_185_[24] ),
    .B(_03612_),
    .Y(_03640_));
 sky130_fd_sc_hd__inv_2 _09231_ (.A(_03613_),
    .Y(_03641_));
 sky130_fd_sc_hd__nand2_1 _09232_ (.A(_02383_),
    .B(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__xnor2_1 _09233_ (.A(_02817_),
    .B(_02787_),
    .Y(_03643_));
 sky130_fd_sc_hd__xnor2_1 _09234_ (.A(_02858_),
    .B(_03643_),
    .Y(_03644_));
 sky130_fd_sc_hd__xnor2_1 _09235_ (.A(\_185_[25] ),
    .B(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__xor2_1 _09236_ (.A(_02422_),
    .B(_03645_),
    .X(_03646_));
 sky130_fd_sc_hd__a21o_1 _09237_ (.A1(_03640_),
    .A2(_03642_),
    .B1(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__nand3_1 _09238_ (.A(_03640_),
    .B(_03642_),
    .C(_03646_),
    .Y(_03648_));
 sky130_fd_sc_hd__and2_1 _09239_ (.A(_03647_),
    .B(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__xnor2_1 _09240_ (.A(_02431_),
    .B(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__a21oi_1 _09241_ (.A1(_03615_),
    .A2(_03619_),
    .B1(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__and3_1 _09242_ (.A(_03615_),
    .B(_03619_),
    .C(_03650_),
    .X(_03652_));
 sky130_fd_sc_hd__or2_1 _09243_ (.A(_03651_),
    .B(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__a21o_1 _09244_ (.A1(\_228_[25] ),
    .A2(\_231_[25] ),
    .B1(_02852_),
    .X(_03654_));
 sky130_fd_sc_hd__o21a_1 _09245_ (.A1(\_228_[25] ),
    .A2(\_231_[25] ),
    .B1(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__xnor2_1 _09246_ (.A(_03653_),
    .B(_03655_),
    .Y(_03656_));
 sky130_fd_sc_hd__o21ai_1 _09247_ (.A1(_03638_),
    .A2(_03639_),
    .B1(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__or3_1 _09248_ (.A(_03638_),
    .B(_03639_),
    .C(_03656_),
    .X(_03658_));
 sky130_fd_sc_hd__and2_1 _09249_ (.A(_03657_),
    .B(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__or2b_1 _09250_ (.A(_03627_),
    .B_N(_03625_),
    .X(_03660_));
 sky130_fd_sc_hd__a21bo_1 _09251_ (.A1(_03628_),
    .A2(_03634_),
    .B1_N(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__xor2_1 _09252_ (.A(_03659_),
    .B(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__nand2_1 _09253_ (.A(\_170_[25] ),
    .B(_02852_),
    .Y(_03663_));
 sky130_fd_sc_hd__or2_1 _09254_ (.A(\_170_[25] ),
    .B(_02852_),
    .X(_03664_));
 sky130_fd_sc_hd__and2_1 _09255_ (.A(_03663_),
    .B(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__o21a_1 _09256_ (.A1(_03600_),
    .A2(_03606_),
    .B1(_03599_),
    .X(_03666_));
 sky130_fd_sc_hd__xnor2_2 _09257_ (.A(_03665_),
    .B(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__or2_1 _09258_ (.A(_01519_),
    .B(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__o211a_1 _09259_ (.A1(_02380_),
    .A2(_03662_),
    .B1(_03668_),
    .C1(_01439_),
    .X(_03669_));
 sky130_fd_sc_hd__a211o_1 _09260_ (.A1(_02852_),
    .A2(_03032_),
    .B1(_03309_),
    .C1(_03669_),
    .X(_00396_));
 sky130_fd_sc_hd__and2b_1 _09261_ (.A_N(_03653_),
    .B(_03655_),
    .X(_03670_));
 sky130_fd_sc_hd__nand2_1 _09262_ (.A(_02431_),
    .B(_03649_),
    .Y(_03671_));
 sky130_fd_sc_hd__nand2_1 _09263_ (.A(\_185_[25] ),
    .B(_03644_),
    .Y(_03672_));
 sky130_fd_sc_hd__inv_2 _09264_ (.A(_03645_),
    .Y(_03673_));
 sky130_fd_sc_hd__nand2_1 _09265_ (.A(_02422_),
    .B(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__xnor2_1 _09266_ (.A(_02820_),
    .B(_02790_),
    .Y(_03675_));
 sky130_fd_sc_hd__xnor2_1 _09267_ (.A(_02862_),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__xnor2_1 _09268_ (.A(\_185_[26] ),
    .B(_03676_),
    .Y(_03677_));
 sky130_fd_sc_hd__xor2_1 _09269_ (.A(_02451_),
    .B(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__a21o_1 _09270_ (.A1(_03672_),
    .A2(_03674_),
    .B1(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__nand3_1 _09271_ (.A(_03672_),
    .B(_03674_),
    .C(_03678_),
    .Y(_03680_));
 sky130_fd_sc_hd__and2_1 _09272_ (.A(_03679_),
    .B(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__xnor2_1 _09273_ (.A(_02460_),
    .B(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__a21oi_1 _09274_ (.A1(_03647_),
    .A2(_03671_),
    .B1(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__and3_1 _09275_ (.A(_03647_),
    .B(_03671_),
    .C(_03682_),
    .X(_03684_));
 sky130_fd_sc_hd__or2_1 _09276_ (.A(_03683_),
    .B(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__a21o_1 _09277_ (.A1(\_228_[26] ),
    .A2(\_231_[26] ),
    .B1(_02855_),
    .X(_03686_));
 sky130_fd_sc_hd__o21a_1 _09278_ (.A1(\_228_[26] ),
    .A2(\_231_[26] ),
    .B1(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__xnor2_1 _09279_ (.A(_03685_),
    .B(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__o21ai_1 _09280_ (.A1(_03651_),
    .A2(_03670_),
    .B1(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__or3_1 _09281_ (.A(_03651_),
    .B(_03670_),
    .C(_03688_),
    .X(_03690_));
 sky130_fd_sc_hd__and2_1 _09282_ (.A(_03689_),
    .B(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__nand2_1 _09283_ (.A(_03628_),
    .B(_03659_),
    .Y(_03692_));
 sky130_fd_sc_hd__a21o_1 _09284_ (.A1(_03630_),
    .A2(_03633_),
    .B1(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__a21bo_1 _09285_ (.A1(_03660_),
    .A2(_03657_),
    .B1_N(_03658_),
    .X(_03694_));
 sky130_fd_sc_hd__nand2_1 _09286_ (.A(_03693_),
    .B(_03694_),
    .Y(_03695_));
 sky130_fd_sc_hd__nand2_1 _09287_ (.A(_03691_),
    .B(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__or2_1 _09288_ (.A(_03691_),
    .B(_03695_),
    .X(_03697_));
 sky130_fd_sc_hd__or2_1 _09289_ (.A(\_170_[26] ),
    .B(_02855_),
    .X(_03698_));
 sky130_fd_sc_hd__nand2_1 _09290_ (.A(\_170_[26] ),
    .B(_02855_),
    .Y(_03699_));
 sky130_fd_sc_hd__nand2_1 _09291_ (.A(_03698_),
    .B(_03699_),
    .Y(_03700_));
 sky130_fd_sc_hd__nor2_1 _09292_ (.A(_03600_),
    .B(_03606_),
    .Y(_03701_));
 sky130_fd_sc_hd__a21boi_1 _09293_ (.A1(_03599_),
    .A2(_03663_),
    .B1_N(_03664_),
    .Y(_03702_));
 sky130_fd_sc_hd__a21o_1 _09294_ (.A1(_03701_),
    .A2(_03664_),
    .B1(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__xnor2_1 _09295_ (.A(_03700_),
    .B(_03703_),
    .Y(_03704_));
 sky130_fd_sc_hd__a21o_1 _09296_ (.A1(_01427_),
    .A2(_03704_),
    .B1(_02002_),
    .X(_03705_));
 sky130_fd_sc_hd__a31o_1 _09297_ (.A1(_01355_),
    .A2(_03696_),
    .A3(_03697_),
    .B1(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__o211a_1 _09298_ (.A1(_02855_),
    .A2(_01426_),
    .B1(_03379_),
    .C1(_03706_),
    .X(_00397_));
 sky130_fd_sc_hd__and2b_1 _09299_ (.A_N(_03685_),
    .B(_03687_),
    .X(_03707_));
 sky130_fd_sc_hd__nand2_1 _09300_ (.A(_02460_),
    .B(_03681_),
    .Y(_03708_));
 sky130_fd_sc_hd__nand2_1 _09301_ (.A(\_185_[26] ),
    .B(_03676_),
    .Y(_03709_));
 sky130_fd_sc_hd__inv_2 _09302_ (.A(_03677_),
    .Y(_03710_));
 sky130_fd_sc_hd__nand2_1 _09303_ (.A(_02451_),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__xnor2_1 _09304_ (.A(_02823_),
    .B(_02794_),
    .Y(_03712_));
 sky130_fd_sc_hd__xnor2_1 _09305_ (.A(_02865_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__nand2_1 _09306_ (.A(\_185_[27] ),
    .B(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__or2_1 _09307_ (.A(\_185_[27] ),
    .B(_03713_),
    .X(_03715_));
 sky130_fd_sc_hd__nand2_1 _09308_ (.A(_03714_),
    .B(_03715_),
    .Y(_03716_));
 sky130_fd_sc_hd__xor2_1 _09309_ (.A(_02486_),
    .B(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__a21o_1 _09310_ (.A1(_03709_),
    .A2(_03711_),
    .B1(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__nand3_1 _09311_ (.A(_03709_),
    .B(_03711_),
    .C(_03717_),
    .Y(_03719_));
 sky130_fd_sc_hd__and2_1 _09312_ (.A(_03718_),
    .B(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__xnor2_1 _09313_ (.A(_02495_),
    .B(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__a21oi_1 _09314_ (.A1(_03679_),
    .A2(_03708_),
    .B1(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__and3_1 _09315_ (.A(_03679_),
    .B(_03708_),
    .C(_03721_),
    .X(_03723_));
 sky130_fd_sc_hd__or2_1 _09316_ (.A(_03722_),
    .B(_03723_),
    .X(_03724_));
 sky130_fd_sc_hd__a21o_1 _09317_ (.A1(\_228_[27] ),
    .A2(\_231_[27] ),
    .B1(_02858_),
    .X(_03725_));
 sky130_fd_sc_hd__o21a_1 _09318_ (.A1(\_228_[27] ),
    .A2(\_231_[27] ),
    .B1(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__xnor2_1 _09319_ (.A(_03724_),
    .B(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__nor3_1 _09320_ (.A(_03683_),
    .B(_03707_),
    .C(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__o21ai_1 _09321_ (.A1(_03683_),
    .A2(_03707_),
    .B1(_03727_),
    .Y(_03729_));
 sky130_fd_sc_hd__and2b_1 _09322_ (.A_N(_03728_),
    .B(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__a21oi_1 _09323_ (.A1(_03689_),
    .A2(_03696_),
    .B1(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__a31o_1 _09324_ (.A1(_03689_),
    .A2(_03696_),
    .A3(_03730_),
    .B1(_01408_),
    .X(_03732_));
 sky130_fd_sc_hd__xnor2_2 _09325_ (.A(\_170_[27] ),
    .B(_02858_),
    .Y(_03733_));
 sky130_fd_sc_hd__a21bo_1 _09326_ (.A1(_03698_),
    .A2(_03703_),
    .B1_N(_03699_),
    .X(_03734_));
 sky130_fd_sc_hd__xor2_2 _09327_ (.A(_03733_),
    .B(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__nand2_1 _09328_ (.A(_02404_),
    .B(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__o211a_1 _09329_ (.A1(_03731_),
    .A2(_03732_),
    .B1(_03736_),
    .C1(_01439_),
    .X(_03737_));
 sky130_fd_sc_hd__a211o_1 _09330_ (.A1(_02858_),
    .A2(_03032_),
    .B1(_03309_),
    .C1(_03737_),
    .X(_00398_));
 sky130_fd_sc_hd__nand2_1 _09331_ (.A(_03691_),
    .B(_03730_),
    .Y(_03738_));
 sky130_fd_sc_hd__o221a_1 _09332_ (.A1(_03689_),
    .A2(_03728_),
    .B1(_03738_),
    .B2(_03694_),
    .C1(_03729_),
    .X(_03739_));
 sky130_fd_sc_hd__a211o_1 _09333_ (.A1(_03630_),
    .A2(_03633_),
    .B1(_03692_),
    .C1(_03738_),
    .X(_03740_));
 sky130_fd_sc_hd__and2b_1 _09334_ (.A_N(_03724_),
    .B(_03726_),
    .X(_03741_));
 sky130_fd_sc_hd__nand2_1 _09335_ (.A(_02495_),
    .B(_03720_),
    .Y(_03742_));
 sky130_fd_sc_hd__nand3_1 _09336_ (.A(_02486_),
    .B(_03714_),
    .C(_03715_),
    .Y(_03743_));
 sky130_fd_sc_hd__xnor2_1 _09337_ (.A(_02827_),
    .B(_02797_),
    .Y(_03744_));
 sky130_fd_sc_hd__xnor2_1 _09338_ (.A(_02868_),
    .B(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__nand2_1 _09339_ (.A(\_185_[28] ),
    .B(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__or2_1 _09340_ (.A(\_185_[28] ),
    .B(_03745_),
    .X(_03747_));
 sky130_fd_sc_hd__nand2_1 _09341_ (.A(_03746_),
    .B(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__xor2_1 _09342_ (.A(_02506_),
    .B(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__a21o_1 _09343_ (.A1(_03714_),
    .A2(_03743_),
    .B1(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__nand3_1 _09344_ (.A(_03714_),
    .B(_03743_),
    .C(_03749_),
    .Y(_03751_));
 sky130_fd_sc_hd__and2_1 _09345_ (.A(_03750_),
    .B(_03751_),
    .X(_03752_));
 sky130_fd_sc_hd__nand2_1 _09346_ (.A(_02514_),
    .B(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__or2_1 _09347_ (.A(_02514_),
    .B(_03752_),
    .X(_03754_));
 sky130_fd_sc_hd__nand2_1 _09348_ (.A(_03753_),
    .B(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__a21oi_1 _09349_ (.A1(_03718_),
    .A2(_03742_),
    .B1(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__and3_1 _09350_ (.A(_03718_),
    .B(_03742_),
    .C(_03755_),
    .X(_03757_));
 sky130_fd_sc_hd__or2_1 _09351_ (.A(_03756_),
    .B(_03757_),
    .X(_03758_));
 sky130_fd_sc_hd__a21o_1 _09352_ (.A1(\_228_[28] ),
    .A2(\_231_[28] ),
    .B1(_02862_),
    .X(_03759_));
 sky130_fd_sc_hd__o21a_1 _09353_ (.A1(\_228_[28] ),
    .A2(\_231_[28] ),
    .B1(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__xnor2_1 _09354_ (.A(_03758_),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__o21ai_2 _09355_ (.A1(_03722_),
    .A2(_03741_),
    .B1(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__or3_1 _09356_ (.A(_03722_),
    .B(_03741_),
    .C(_03761_),
    .X(_03763_));
 sky130_fd_sc_hd__nand2_1 _09357_ (.A(_03762_),
    .B(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__a21o_1 _09358_ (.A1(_03739_),
    .A2(_03740_),
    .B1(_03764_),
    .X(_03765_));
 sky130_fd_sc_hd__a31oi_1 _09359_ (.A1(_03764_),
    .A2(_03739_),
    .A3(_03740_),
    .B1(_01923_),
    .Y(_03766_));
 sky130_fd_sc_hd__nor2_1 _09360_ (.A(_03700_),
    .B(_03733_),
    .Y(_03767_));
 sky130_fd_sc_hd__o211a_1 _09361_ (.A1(\_170_[27] ),
    .A2(_02858_),
    .B1(_02855_),
    .C1(\_170_[26] ),
    .X(_03768_));
 sky130_fd_sc_hd__a221o_1 _09362_ (.A1(\_170_[27] ),
    .A2(_02858_),
    .B1(_03702_),
    .B2(_03767_),
    .C1(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__a31o_1 _09363_ (.A1(_03701_),
    .A2(_03665_),
    .A3(_03767_),
    .B1(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__or2_1 _09364_ (.A(\_170_[28] ),
    .B(_02862_),
    .X(_03771_));
 sky130_fd_sc_hd__nand2_1 _09365_ (.A(\_170_[28] ),
    .B(_02862_),
    .Y(_03772_));
 sky130_fd_sc_hd__nand2_1 _09366_ (.A(_03771_),
    .B(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__xnor2_1 _09367_ (.A(_03770_),
    .B(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__and2_1 _09368_ (.A(_01437_),
    .B(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__a211o_1 _09369_ (.A1(_03765_),
    .A2(_03766_),
    .B1(_03775_),
    .C1(_01495_),
    .X(_03776_));
 sky130_fd_sc_hd__o211a_1 _09370_ (.A1(_02862_),
    .A2(_01426_),
    .B1(_03379_),
    .C1(_03776_),
    .X(_00399_));
 sky130_fd_sc_hd__and2b_1 _09371_ (.A_N(_03758_),
    .B(_03760_),
    .X(_03777_));
 sky130_fd_sc_hd__nand3_1 _09372_ (.A(_02506_),
    .B(_03746_),
    .C(_03747_),
    .Y(_03778_));
 sky130_fd_sc_hd__xnor2_1 _09373_ (.A(_02830_),
    .B(_02801_),
    .Y(_03779_));
 sky130_fd_sc_hd__xnor2_1 _09374_ (.A(_02871_),
    .B(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__nand2_1 _09375_ (.A(\_185_[29] ),
    .B(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__or2_1 _09376_ (.A(\_185_[29] ),
    .B(_03780_),
    .X(_03782_));
 sky130_fd_sc_hd__nand2_1 _09377_ (.A(_03781_),
    .B(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__inv_2 _09378_ (.A(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__nand2_1 _09379_ (.A(_02540_),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__or2_1 _09380_ (.A(_02540_),
    .B(_03784_),
    .X(_03786_));
 sky130_fd_sc_hd__nand2_1 _09381_ (.A(_03785_),
    .B(_03786_),
    .Y(_03787_));
 sky130_fd_sc_hd__a21o_1 _09382_ (.A1(_03746_),
    .A2(_03778_),
    .B1(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__nand3_1 _09383_ (.A(_03746_),
    .B(_03778_),
    .C(_03787_),
    .Y(_03789_));
 sky130_fd_sc_hd__and2_1 _09384_ (.A(_03788_),
    .B(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__nand2_1 _09385_ (.A(_02549_),
    .B(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__or2_1 _09386_ (.A(_02549_),
    .B(_03790_),
    .X(_03792_));
 sky130_fd_sc_hd__nand2_1 _09387_ (.A(_03791_),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__a21oi_1 _09388_ (.A1(_03750_),
    .A2(_03753_),
    .B1(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__and3_1 _09389_ (.A(_03750_),
    .B(_03753_),
    .C(_03793_),
    .X(_03795_));
 sky130_fd_sc_hd__or2_1 _09390_ (.A(_03794_),
    .B(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__a21o_1 _09391_ (.A1(\_228_[29] ),
    .A2(\_231_[29] ),
    .B1(_02865_),
    .X(_03797_));
 sky130_fd_sc_hd__o21a_1 _09392_ (.A1(\_228_[29] ),
    .A2(\_231_[29] ),
    .B1(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__xnor2_1 _09393_ (.A(_03796_),
    .B(_03798_),
    .Y(_03799_));
 sky130_fd_sc_hd__o21ai_1 _09394_ (.A1(_03756_),
    .A2(_03777_),
    .B1(_03799_),
    .Y(_03800_));
 sky130_fd_sc_hd__inv_2 _09395_ (.A(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__nor3_1 _09396_ (.A(_03756_),
    .B(_03777_),
    .C(_03799_),
    .Y(_03802_));
 sky130_fd_sc_hd__nor2_1 _09397_ (.A(_03801_),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__and3_1 _09398_ (.A(_03762_),
    .B(_03765_),
    .C(_03803_),
    .X(_03804_));
 sky130_fd_sc_hd__a21oi_1 _09399_ (.A1(_03762_),
    .A2(_03765_),
    .B1(_03803_),
    .Y(_03805_));
 sky130_fd_sc_hd__or2_1 _09400_ (.A(\_170_[29] ),
    .B(_02865_),
    .X(_03806_));
 sky130_fd_sc_hd__nand2_1 _09401_ (.A(\_170_[29] ),
    .B(_02865_),
    .Y(_03807_));
 sky130_fd_sc_hd__nand2_1 _09402_ (.A(_03806_),
    .B(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__a21bo_1 _09403_ (.A1(_03770_),
    .A2(_03771_),
    .B1_N(_03772_),
    .X(_03809_));
 sky130_fd_sc_hd__xnor2_2 _09404_ (.A(_03808_),
    .B(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__or2_1 _09405_ (.A(_01519_),
    .B(_03810_),
    .X(_03811_));
 sky130_fd_sc_hd__o311a_1 _09406_ (.A1(_01409_),
    .A2(_03804_),
    .A3(_03805_),
    .B1(_03811_),
    .C1(_01799_),
    .X(_03812_));
 sky130_fd_sc_hd__a211o_1 _09407_ (.A1(_02865_),
    .A2(_01884_),
    .B1(_03309_),
    .C1(_03812_),
    .X(_00400_));
 sky130_fd_sc_hd__and2b_1 _09408_ (.A_N(_03796_),
    .B(_03798_),
    .X(_03813_));
 sky130_fd_sc_hd__inv_2 _09409_ (.A(_02573_),
    .Y(_03814_));
 sky130_fd_sc_hd__xnor2_1 _09410_ (.A(_02804_),
    .B(_02768_),
    .Y(_03815_));
 sky130_fd_sc_hd__xnor2_1 _09411_ (.A(_02835_),
    .B(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__nand2_1 _09412_ (.A(\_185_[30] ),
    .B(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__or2_1 _09413_ (.A(\_185_[30] ),
    .B(_03816_),
    .X(_03818_));
 sky130_fd_sc_hd__nand2_1 _09414_ (.A(_03817_),
    .B(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__xnor2_1 _09415_ (.A(_03814_),
    .B(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__a21oi_1 _09416_ (.A1(_03781_),
    .A2(_03785_),
    .B1(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__and3_1 _09417_ (.A(_03781_),
    .B(_03785_),
    .C(_03820_),
    .X(_03822_));
 sky130_fd_sc_hd__nor2_1 _09418_ (.A(_03821_),
    .B(_03822_),
    .Y(_03823_));
 sky130_fd_sc_hd__xnor2_1 _09419_ (.A(_02582_),
    .B(_03823_),
    .Y(_03824_));
 sky130_fd_sc_hd__a21o_1 _09420_ (.A1(_03788_),
    .A2(_03791_),
    .B1(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__nand3_1 _09421_ (.A(_03788_),
    .B(_03791_),
    .C(_03824_),
    .Y(_03826_));
 sky130_fd_sc_hd__a21o_1 _09422_ (.A1(\_228_[30] ),
    .A2(\_231_[30] ),
    .B1(_02868_),
    .X(_03827_));
 sky130_fd_sc_hd__o21a_1 _09423_ (.A1(\_228_[30] ),
    .A2(\_231_[30] ),
    .B1(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__and3_1 _09424_ (.A(_03825_),
    .B(_03826_),
    .C(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__a21oi_1 _09425_ (.A1(_03825_),
    .A2(_03826_),
    .B1(_03828_),
    .Y(_03830_));
 sky130_fd_sc_hd__nor2_1 _09426_ (.A(_03829_),
    .B(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__o21ai_1 _09427_ (.A1(_03794_),
    .A2(_03813_),
    .B1(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__or3_1 _09428_ (.A(_03794_),
    .B(_03813_),
    .C(_03831_),
    .X(_03833_));
 sky130_fd_sc_hd__nand2_1 _09429_ (.A(_03832_),
    .B(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__a31o_1 _09430_ (.A1(_03762_),
    .A2(_03765_),
    .A3(_03800_),
    .B1(_03802_),
    .X(_03835_));
 sky130_fd_sc_hd__xor2_1 _09431_ (.A(_03834_),
    .B(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__nand2_1 _09432_ (.A(\_170_[30] ),
    .B(_02868_),
    .Y(_03837_));
 sky130_fd_sc_hd__or2_1 _09433_ (.A(\_170_[30] ),
    .B(_02868_),
    .X(_03838_));
 sky130_fd_sc_hd__nand2_1 _09434_ (.A(_03837_),
    .B(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__a21bo_1 _09435_ (.A1(_03806_),
    .A2(_03809_),
    .B1_N(_03807_),
    .X(_03840_));
 sky130_fd_sc_hd__xor2_2 _09436_ (.A(_03839_),
    .B(_03840_),
    .X(_03841_));
 sky130_fd_sc_hd__nand2_1 _09437_ (.A(_02404_),
    .B(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__o211a_1 _09438_ (.A1(_02380_),
    .A2(_03836_),
    .B1(_03842_),
    .C1(_01439_),
    .X(_03843_));
 sky130_fd_sc_hd__a211o_1 _09439_ (.A1(_02868_),
    .A2(_01884_),
    .B1(_03309_),
    .C1(_03843_),
    .X(_00401_));
 sky130_fd_sc_hd__a311o_1 _09440_ (.A1(_03762_),
    .A2(_03765_),
    .A3(_03800_),
    .B1(_03802_),
    .C1(_03834_),
    .X(_03844_));
 sky130_fd_sc_hd__a21bo_1 _09441_ (.A1(_03826_),
    .A2(_03828_),
    .B1_N(_03825_),
    .X(_03845_));
 sky130_fd_sc_hd__a21oi_1 _09442_ (.A1(_02582_),
    .A2(_03823_),
    .B1(_03821_),
    .Y(_03846_));
 sky130_fd_sc_hd__xnor2_1 _09443_ (.A(_02807_),
    .B(_02772_),
    .Y(_03847_));
 sky130_fd_sc_hd__a21o_1 _09444_ (.A1(_02871_),
    .A2(\_231_[31] ),
    .B1(\_228_[31] ),
    .X(_03848_));
 sky130_fd_sc_hd__o21a_1 _09445_ (.A1(_02871_),
    .A2(\_231_[31] ),
    .B1(_03848_),
    .X(_03849_));
 sky130_fd_sc_hd__xnor2_1 _09446_ (.A(_03847_),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__xnor2_1 _09447_ (.A(_02598_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__o21ai_1 _09448_ (.A1(_03814_),
    .A2(_03819_),
    .B1(_03817_),
    .Y(_03852_));
 sky130_fd_sc_hd__xnor2_1 _09449_ (.A(_02839_),
    .B(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hd__xnor2_1 _09450_ (.A(_03851_),
    .B(_03853_),
    .Y(_03854_));
 sky130_fd_sc_hd__xnor2_1 _09451_ (.A(_03846_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__xnor2_1 _09452_ (.A(_03845_),
    .B(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__and3_1 _09453_ (.A(_03832_),
    .B(_03844_),
    .C(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__a21oi_1 _09454_ (.A1(_03832_),
    .A2(_03844_),
    .B1(_03856_),
    .Y(_03858_));
 sky130_fd_sc_hd__or3_1 _09455_ (.A(_01923_),
    .B(_03857_),
    .C(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__a21bo_1 _09456_ (.A1(_03838_),
    .A2(_03840_),
    .B1_N(_03837_),
    .X(_03860_));
 sky130_fd_sc_hd__xnor2_1 _09457_ (.A(\_170_[31] ),
    .B(_02871_),
    .Y(_03861_));
 sky130_fd_sc_hd__xnor2_2 _09458_ (.A(_03860_),
    .B(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__a21oi_1 _09459_ (.A1(_01856_),
    .A2(_03862_),
    .B1(_01884_),
    .Y(_03863_));
 sky130_fd_sc_hd__buf_6 _09460_ (.A(_01423_),
    .X(_03864_));
 sky130_fd_sc_hd__o21ai_1 _09461_ (.A1(_02871_),
    .A2(_01421_),
    .B1(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__a21oi_1 _09462_ (.A1(_03859_),
    .A2(_03863_),
    .B1(_03865_),
    .Y(_00402_));
 sky130_fd_sc_hd__buf_6 _09463_ (.A(_01418_),
    .X(_03866_));
 sky130_fd_sc_hd__inv_2 _09464_ (.A(_03866_),
    .Y(_00106_));
 sky130_fd_sc_hd__inv_2 _09465_ (.A(_03866_),
    .Y(_00107_));
 sky130_fd_sc_hd__inv_2 _09466_ (.A(_03866_),
    .Y(_00108_));
 sky130_fd_sc_hd__inv_2 _09467_ (.A(_03866_),
    .Y(_00109_));
 sky130_fd_sc_hd__inv_2 _09468_ (.A(_03866_),
    .Y(_00110_));
 sky130_fd_sc_hd__o211ai_4 _09469_ (.A1(_01295_),
    .A2(_01271_),
    .B1(_01272_),
    .C1(_01274_),
    .Y(_03867_));
 sky130_fd_sc_hd__clkbuf_4 _09470_ (.A(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__buf_2 _09471_ (.A(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__clkbuf_4 _09472_ (.A(_03867_),
    .X(_03870_));
 sky130_fd_sc_hd__clkbuf_4 _09473_ (.A(_01230_),
    .X(_03871_));
 sky130_fd_sc_hd__buf_2 _09474_ (.A(_01234_),
    .X(_03872_));
 sky130_fd_sc_hd__nand2b_4 _09475_ (.A_N(_01280_),
    .B(_01283_),
    .Y(_03873_));
 sky130_fd_sc_hd__buf_2 _09476_ (.A(\_195_[2] ),
    .X(_03874_));
 sky130_fd_sc_hd__nor2_4 _09477_ (.A(_03874_),
    .B(_01282_),
    .Y(_03875_));
 sky130_fd_sc_hd__nor2_4 _09478_ (.A(\_195_[3] ),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__xor2_1 _09479_ (.A(\_195_[1] ),
    .B(\_195_[0] ),
    .X(_03877_));
 sky130_fd_sc_hd__buf_4 _09480_ (.A(_03877_),
    .X(_03878_));
 sky130_fd_sc_hd__clkinv_2 _09481_ (.A(\_195_[3] ),
    .Y(_03879_));
 sky130_fd_sc_hd__nor2_4 _09482_ (.A(_03879_),
    .B(_03875_),
    .Y(_03880_));
 sky130_fd_sc_hd__a22o_1 _09483_ (.A1(_03873_),
    .A2(_03876_),
    .B1(_03878_),
    .B2(_03880_),
    .X(_03881_));
 sky130_fd_sc_hd__nand2_1 _09484_ (.A(_03872_),
    .B(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__or2_1 _09485_ (.A(_01277_),
    .B(_03878_),
    .X(_03883_));
 sky130_fd_sc_hd__buf_2 _09486_ (.A(_01240_),
    .X(_03884_));
 sky130_fd_sc_hd__and2_1 _09487_ (.A(_01277_),
    .B(_01282_),
    .X(_03885_));
 sky130_fd_sc_hd__buf_2 _09488_ (.A(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__nor2_1 _09489_ (.A(_03884_),
    .B(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__nand2b_4 _09490_ (.A_N(_01282_),
    .B(_01278_),
    .Y(_03888_));
 sky130_fd_sc_hd__or2_1 _09491_ (.A(\_195_[2] ),
    .B(\_195_[1] ),
    .X(_03889_));
 sky130_fd_sc_hd__clkbuf_4 _09492_ (.A(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__or2b_1 _09493_ (.A(_03874_),
    .B_N(\_195_[0] ),
    .X(_03891_));
 sky130_fd_sc_hd__and3_1 _09494_ (.A(_01240_),
    .B(_03890_),
    .C(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__buf_2 _09495_ (.A(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__a21o_1 _09496_ (.A1(_03888_),
    .A2(_03893_),
    .B1(_01234_),
    .X(_03894_));
 sky130_fd_sc_hd__a21o_1 _09497_ (.A1(_03883_),
    .A2(_03887_),
    .B1(_03894_),
    .X(_03895_));
 sky130_fd_sc_hd__clkbuf_4 _09498_ (.A(_03891_),
    .X(_03896_));
 sky130_fd_sc_hd__nor2b_4 _09499_ (.A(_01282_),
    .B_N(_03874_),
    .Y(_03897_));
 sky130_fd_sc_hd__nand2_2 _09500_ (.A(_01280_),
    .B(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__and3_1 _09501_ (.A(_01241_),
    .B(_03896_),
    .C(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__or2b_1 _09502_ (.A(_01279_),
    .B_N(_03874_),
    .X(_03900_));
 sky130_fd_sc_hd__clkbuf_4 _09503_ (.A(_03900_),
    .X(_03901_));
 sky130_fd_sc_hd__or2b_1 _09504_ (.A(_03874_),
    .B_N(_01279_),
    .X(_03902_));
 sky130_fd_sc_hd__clkbuf_4 _09505_ (.A(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__nand2_1 _09506_ (.A(_03901_),
    .B(_03903_),
    .Y(_03904_));
 sky130_fd_sc_hd__or2_1 _09507_ (.A(_01240_),
    .B(_01283_),
    .X(_03905_));
 sky130_fd_sc_hd__nor2_1 _09508_ (.A(_03904_),
    .B(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__or2_2 _09509_ (.A(_01240_),
    .B(_01280_),
    .X(_03907_));
 sky130_fd_sc_hd__nor2_1 _09510_ (.A(_01283_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__o21ai_1 _09511_ (.A1(_03880_),
    .A2(_03908_),
    .B1(_01235_),
    .Y(_03909_));
 sky130_fd_sc_hd__inv_2 _09512_ (.A(\_195_[5] ),
    .Y(_03910_));
 sky130_fd_sc_hd__o311a_1 _09513_ (.A1(_01235_),
    .A2(_03899_),
    .A3(_03906_),
    .B1(_03909_),
    .C1(_03910_),
    .X(_03911_));
 sky130_fd_sc_hd__a31o_1 _09514_ (.A1(_03871_),
    .A2(_03882_),
    .A3(_03895_),
    .B1(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__o32ai_4 _09515_ (.A1(\_392_[4] ),
    .A2(_01206_),
    .A3(_01246_),
    .B1(_01268_),
    .B2(_01251_),
    .Y(_03913_));
 sky130_fd_sc_hd__buf_2 _09516_ (.A(_03913_),
    .X(_03914_));
 sky130_fd_sc_hd__o221a_2 _09517_ (.A1(\_246_[0] ),
    .A2(_01314_),
    .B1(_03914_),
    .B2(\_243_[0] ),
    .C1(_01413_),
    .X(_03915_));
 sky130_fd_sc_hd__xnor2_1 _09518_ (.A(\_142_[0] ),
    .B(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__xnor2_1 _09519_ (.A(_03912_),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__nand2_1 _09520_ (.A(_03870_),
    .B(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__o211a_1 _09521_ (.A1(\_185_[0] ),
    .A2(_03869_),
    .B1(_03379_),
    .C1(_03918_),
    .X(_00409_));
 sky130_fd_sc_hd__buf_2 _09522_ (.A(_02833_),
    .X(_03919_));
 sky130_fd_sc_hd__o2bb2ai_1 _09523_ (.A1_N(\_142_[0] ),
    .A2_N(_03915_),
    .B1(_03916_),
    .B2(_03912_),
    .Y(_03920_));
 sky130_fd_sc_hd__o221a_1 _09524_ (.A1(\_246_[1] ),
    .A2(_01313_),
    .B1(_03913_),
    .B2(\_243_[1] ),
    .C1(_01429_),
    .X(_03921_));
 sky130_fd_sc_hd__xor2_1 _09525_ (.A(\_142_[1] ),
    .B(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__nor2_1 _09526_ (.A(\_195_[1] ),
    .B(\_195_[0] ),
    .Y(_03923_));
 sky130_fd_sc_hd__or3_1 _09527_ (.A(_03874_),
    .B(_01291_),
    .C(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__buf_2 _09528_ (.A(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__mux2_1 _09529_ (.A0(_03883_),
    .A1(_03925_),
    .S(_01240_),
    .X(_03926_));
 sky130_fd_sc_hd__nand2_4 _09530_ (.A(_01277_),
    .B(_03878_),
    .Y(_03927_));
 sky130_fd_sc_hd__or3b_4 _09531_ (.A(_01279_),
    .B(\_195_[0] ),
    .C_N(_03874_),
    .X(_03928_));
 sky130_fd_sc_hd__or3b_2 _09532_ (.A(_03874_),
    .B(\_195_[0] ),
    .C_N(_01279_),
    .X(_03929_));
 sky130_fd_sc_hd__a31o_1 _09533_ (.A1(_03879_),
    .A2(_03928_),
    .A3(_03929_),
    .B1(\_195_[4] ),
    .X(_03930_));
 sky130_fd_sc_hd__a31oi_1 _09534_ (.A1(_01241_),
    .A2(_03903_),
    .A3(_03927_),
    .B1(_03930_),
    .Y(_03931_));
 sky130_fd_sc_hd__a31o_1 _09535_ (.A1(_01234_),
    .A2(_03898_),
    .A3(_03926_),
    .B1(_03931_),
    .X(_03932_));
 sky130_fd_sc_hd__clkinv_2 _09536_ (.A(_01234_),
    .Y(_03933_));
 sky130_fd_sc_hd__nand2_1 _09537_ (.A(_01241_),
    .B(_03896_),
    .Y(_03934_));
 sky130_fd_sc_hd__and3b_2 _09538_ (.A_N(_01277_),
    .B(_01279_),
    .C(_01282_),
    .X(_03935_));
 sky130_fd_sc_hd__and2_1 _09539_ (.A(_01277_),
    .B(_03877_),
    .X(_03936_));
 sky130_fd_sc_hd__or3_1 _09540_ (.A(_01240_),
    .B(_03935_),
    .C(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__or3b_2 _09541_ (.A(\_195_[3] ),
    .B(_03874_),
    .C_N(\_195_[0] ),
    .X(_03938_));
 sky130_fd_sc_hd__a31o_1 _09542_ (.A1(_01234_),
    .A2(_03903_),
    .A3(_03938_),
    .B1(_03910_),
    .X(_03939_));
 sky130_fd_sc_hd__a31o_1 _09543_ (.A1(_03933_),
    .A2(_03934_),
    .A3(_03937_),
    .B1(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__o21ai_1 _09544_ (.A1(_03871_),
    .A2(_03932_),
    .B1(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__xnor2_1 _09545_ (.A(_03922_),
    .B(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__nand2_1 _09546_ (.A(_03920_),
    .B(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__or2_1 _09547_ (.A(_03920_),
    .B(_03942_),
    .X(_03944_));
 sky130_fd_sc_hd__clkbuf_4 _09548_ (.A(_01275_),
    .X(_03945_));
 sky130_fd_sc_hd__buf_2 _09549_ (.A(_03945_),
    .X(_03946_));
 sky130_fd_sc_hd__a21o_1 _09550_ (.A1(_03943_),
    .A2(_03944_),
    .B1(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__o211a_1 _09551_ (.A1(\_185_[1] ),
    .A2(_03869_),
    .B1(_03919_),
    .C1(_03947_),
    .X(_00410_));
 sky130_fd_sc_hd__and2_1 _09552_ (.A(\_142_[1] ),
    .B(_03921_),
    .X(_03948_));
 sky130_fd_sc_hd__o211a_1 _09553_ (.A1(_01230_),
    .A2(_03932_),
    .B1(_03940_),
    .C1(_03922_),
    .X(_03949_));
 sky130_fd_sc_hd__nand2_2 _09554_ (.A(\_195_[2] ),
    .B(\_195_[1] ),
    .Y(_03950_));
 sky130_fd_sc_hd__and2_1 _09555_ (.A(_03879_),
    .B(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__buf_2 _09556_ (.A(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__a221o_1 _09557_ (.A1(_01240_),
    .A2(_03927_),
    .B1(_03952_),
    .B2(_01283_),
    .C1(\_195_[4] ),
    .X(_03953_));
 sky130_fd_sc_hd__nand2_1 _09558_ (.A(_01280_),
    .B(_01282_),
    .Y(_03954_));
 sky130_fd_sc_hd__a32o_1 _09559_ (.A1(_03954_),
    .A2(_03901_),
    .A3(_03938_),
    .B1(_03935_),
    .B2(_03879_),
    .X(_03955_));
 sky130_fd_sc_hd__nand2_1 _09560_ (.A(_01234_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__or2b_1 _09561_ (.A(_01282_),
    .B_N(_01279_),
    .X(_03957_));
 sky130_fd_sc_hd__and2b_1 _09562_ (.A_N(_01277_),
    .B(\_195_[3] ),
    .X(_03958_));
 sky130_fd_sc_hd__a21oi_1 _09563_ (.A1(_03957_),
    .A2(_03958_),
    .B1(\_195_[4] ),
    .Y(_03959_));
 sky130_fd_sc_hd__nand2_2 _09564_ (.A(_01277_),
    .B(_01282_),
    .Y(_03960_));
 sky130_fd_sc_hd__o21ba_1 _09565_ (.A1(_01277_),
    .A2(_01279_),
    .B1_N(\_195_[3] ),
    .X(_03961_));
 sky130_fd_sc_hd__o221a_1 _09566_ (.A1(_01240_),
    .A2(_03960_),
    .B1(_03961_),
    .B2(_01282_),
    .C1(\_195_[4] ),
    .X(_03962_));
 sky130_fd_sc_hd__a211oi_1 _09567_ (.A1(_03907_),
    .A2(_03959_),
    .B1(_03962_),
    .C1(\_195_[5] ),
    .Y(_03963_));
 sky130_fd_sc_hd__a31o_1 _09568_ (.A1(\_195_[5] ),
    .A2(_03953_),
    .A3(_03956_),
    .B1(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__o221a_1 _09569_ (.A1(\_246_[2] ),
    .A2(_01313_),
    .B1(_03913_),
    .B2(\_243_[2] ),
    .C1(_01432_),
    .X(_03965_));
 sky130_fd_sc_hd__xnor2_1 _09570_ (.A(\_142_[2] ),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__xor2_1 _09571_ (.A(_03964_),
    .B(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__o21a_1 _09572_ (.A1(_03948_),
    .A2(_03949_),
    .B1(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__nor3_1 _09573_ (.A(_03948_),
    .B(_03949_),
    .C(_03967_),
    .Y(_03969_));
 sky130_fd_sc_hd__or3_1 _09574_ (.A(_03943_),
    .B(_03968_),
    .C(_03969_),
    .X(_03970_));
 sky130_fd_sc_hd__o21ai_1 _09575_ (.A1(_03968_),
    .A2(_03969_),
    .B1(_03943_),
    .Y(_03971_));
 sky130_fd_sc_hd__a21o_1 _09576_ (.A1(_03970_),
    .A2(_03971_),
    .B1(_03946_),
    .X(_03972_));
 sky130_fd_sc_hd__o211a_1 _09577_ (.A1(\_185_[2] ),
    .A2(_03869_),
    .B1(_03919_),
    .C1(_03972_),
    .X(_00411_));
 sky130_fd_sc_hd__o2bb2ai_1 _09578_ (.A1_N(\_142_[2] ),
    .A2_N(_03965_),
    .B1(_03966_),
    .B2(_03964_),
    .Y(_03973_));
 sky130_fd_sc_hd__o221a_2 _09579_ (.A1(\_246_[3] ),
    .A2(_01313_),
    .B1(_03914_),
    .B2(\_243_[3] ),
    .C1(_01440_),
    .X(_03974_));
 sky130_fd_sc_hd__xnor2_1 _09580_ (.A(\_142_[3] ),
    .B(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__nor2_2 _09581_ (.A(_01278_),
    .B(_03873_),
    .Y(_03976_));
 sky130_fd_sc_hd__nand2_1 _09582_ (.A(_01241_),
    .B(_03888_),
    .Y(_03977_));
 sky130_fd_sc_hd__nor3_1 _09583_ (.A(_01235_),
    .B(_03976_),
    .C(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__nor2_2 _09584_ (.A(_01241_),
    .B(_03878_),
    .Y(_03979_));
 sky130_fd_sc_hd__a211o_1 _09585_ (.A1(_03901_),
    .A2(_03893_),
    .B1(_03979_),
    .C1(_03910_),
    .X(_03980_));
 sky130_fd_sc_hd__nand2_1 _09586_ (.A(_01241_),
    .B(_03925_),
    .Y(_03981_));
 sky130_fd_sc_hd__o31a_1 _09587_ (.A1(_01240_),
    .A2(_01278_),
    .A3(_01291_),
    .B1(_01234_),
    .X(_03982_));
 sky130_fd_sc_hd__nor2b_4 _09588_ (.A(_01279_),
    .B_N(_03874_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_4 _09589_ (.A(_01283_),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__a221o_1 _09590_ (.A1(_03876_),
    .A2(_03928_),
    .B1(_03984_),
    .B2(_03880_),
    .C1(\_195_[4] ),
    .X(_03985_));
 sky130_fd_sc_hd__a21bo_1 _09591_ (.A1(_03981_),
    .A2(_03982_),
    .B1_N(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__a2bb2o_1 _09592_ (.A1_N(_03978_),
    .A2_N(_03980_),
    .B1(_03986_),
    .B2(_03910_),
    .X(_03987_));
 sky130_fd_sc_hd__xor2_1 _09593_ (.A(_03975_),
    .B(_03987_),
    .X(_03988_));
 sky130_fd_sc_hd__xnor2_1 _09594_ (.A(_03973_),
    .B(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__or3_1 _09595_ (.A(_03948_),
    .B(_03949_),
    .C(_03967_),
    .X(_03990_));
 sky130_fd_sc_hd__a31o_1 _09596_ (.A1(_03920_),
    .A2(_03942_),
    .A3(_03990_),
    .B1(_03968_),
    .X(_03991_));
 sky130_fd_sc_hd__nand2_1 _09597_ (.A(_03989_),
    .B(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__or2_1 _09598_ (.A(_03989_),
    .B(_03991_),
    .X(_03993_));
 sky130_fd_sc_hd__a21o_1 _09599_ (.A1(_03992_),
    .A2(_03993_),
    .B1(_03946_),
    .X(_03994_));
 sky130_fd_sc_hd__o211a_1 _09600_ (.A1(\_185_[3] ),
    .A2(_03869_),
    .B1(_03919_),
    .C1(_03994_),
    .X(_00412_));
 sky130_fd_sc_hd__and2b_1 _09601_ (.A_N(_03988_),
    .B(_03973_),
    .X(_03995_));
 sky130_fd_sc_hd__a21oi_1 _09602_ (.A1(_03989_),
    .A2(_03991_),
    .B1(_03995_),
    .Y(_03996_));
 sky130_fd_sc_hd__o221a_1 _09603_ (.A1(\_246_[4] ),
    .A2(_01313_),
    .B1(_03913_),
    .B2(\_243_[4] ),
    .C1(_01442_),
    .X(_03997_));
 sky130_fd_sc_hd__and2_1 _09604_ (.A(\_142_[4] ),
    .B(_03997_),
    .X(_03998_));
 sky130_fd_sc_hd__nor2_1 _09605_ (.A(\_142_[4] ),
    .B(_03997_),
    .Y(_03999_));
 sky130_fd_sc_hd__or2_1 _09606_ (.A(_03998_),
    .B(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__a21oi_1 _09607_ (.A1(_03873_),
    .A2(_03893_),
    .B1(_03979_),
    .Y(_04001_));
 sky130_fd_sc_hd__buf_2 _09608_ (.A(_03879_),
    .X(_04002_));
 sky130_fd_sc_hd__a31oi_1 _09609_ (.A1(_03890_),
    .A2(_03896_),
    .A3(_03927_),
    .B1(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__and2b_1 _09610_ (.A_N(_01277_),
    .B(_01279_),
    .X(_04004_));
 sky130_fd_sc_hd__buf_2 _09611_ (.A(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__nor2_2 _09612_ (.A(_01241_),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__a31o_1 _09613_ (.A1(_03901_),
    .A2(_04006_),
    .A3(_03873_),
    .B1(_01234_),
    .X(_04007_));
 sky130_fd_sc_hd__o221a_1 _09614_ (.A1(_03933_),
    .A2(_04001_),
    .B1(_04003_),
    .B2(_04007_),
    .C1(_01230_),
    .X(_04008_));
 sky130_fd_sc_hd__a311o_1 _09615_ (.A1(_04002_),
    .A2(_03957_),
    .A3(_03903_),
    .B1(_03899_),
    .C1(_01235_),
    .X(_04009_));
 sky130_fd_sc_hd__nor2b_4 _09616_ (.A(_01280_),
    .B_N(_03875_),
    .Y(_04010_));
 sky130_fd_sc_hd__nor2_1 _09617_ (.A(_04010_),
    .B(_03977_),
    .Y(_04011_));
 sky130_fd_sc_hd__o21ai_1 _09618_ (.A1(_03952_),
    .A2(_04011_),
    .B1(_03872_),
    .Y(_04012_));
 sky130_fd_sc_hd__a21oi_1 _09619_ (.A1(_04009_),
    .A2(_04012_),
    .B1(_03871_),
    .Y(_04013_));
 sky130_fd_sc_hd__or2_1 _09620_ (.A(_04008_),
    .B(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__xnor2_1 _09621_ (.A(_04000_),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__or2b_1 _09622_ (.A(_03975_),
    .B_N(_03987_),
    .X(_04016_));
 sky130_fd_sc_hd__a21bo_1 _09623_ (.A1(\_142_[3] ),
    .A2(_03974_),
    .B1_N(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__xor2_2 _09624_ (.A(_04015_),
    .B(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__or2_1 _09625_ (.A(_03996_),
    .B(_04018_),
    .X(_04019_));
 sky130_fd_sc_hd__nand2_1 _09626_ (.A(_03996_),
    .B(_04018_),
    .Y(_04020_));
 sky130_fd_sc_hd__a21o_1 _09627_ (.A1(_04019_),
    .A2(_04020_),
    .B1(_03946_),
    .X(_04021_));
 sky130_fd_sc_hd__o211a_1 _09628_ (.A1(\_185_[4] ),
    .A2(_03869_),
    .B1(_03919_),
    .C1(_04021_),
    .X(_00413_));
 sky130_fd_sc_hd__nor2_1 _09629_ (.A(_04000_),
    .B(_04014_),
    .Y(_04022_));
 sky130_fd_sc_hd__o221a_1 _09630_ (.A1(\_246_[5] ),
    .A2(_01313_),
    .B1(_03914_),
    .B2(\_243_[5] ),
    .C1(_01445_),
    .X(_04023_));
 sky130_fd_sc_hd__xnor2_1 _09631_ (.A(\_142_[5] ),
    .B(_04023_),
    .Y(_04024_));
 sky130_fd_sc_hd__nand2_1 _09632_ (.A(_03903_),
    .B(_03880_),
    .Y(_04025_));
 sky130_fd_sc_hd__nor2_1 _09633_ (.A(_03886_),
    .B(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__nor2_1 _09634_ (.A(_01280_),
    .B(_03888_),
    .Y(_04027_));
 sky130_fd_sc_hd__a21oi_1 _09635_ (.A1(_03884_),
    .A2(_04005_),
    .B1(_03933_),
    .Y(_04028_));
 sky130_fd_sc_hd__o31ai_1 _09636_ (.A1(_03884_),
    .A2(_01292_),
    .A3(_04027_),
    .B1(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__o311a_1 _09637_ (.A1(_01235_),
    .A2(_03979_),
    .A3(_04026_),
    .B1(_04029_),
    .C1(_01230_),
    .X(_04030_));
 sky130_fd_sc_hd__o21ai_1 _09638_ (.A1(_01280_),
    .A2(_03896_),
    .B1(_03950_),
    .Y(_04031_));
 sky130_fd_sc_hd__nor2_1 _09639_ (.A(_03977_),
    .B(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__a211oi_1 _09640_ (.A1(_03901_),
    .A2(_03977_),
    .B1(_04032_),
    .C1(_03933_),
    .Y(_04033_));
 sky130_fd_sc_hd__a211oi_1 _09641_ (.A1(_03937_),
    .A2(_03959_),
    .B1(_04033_),
    .C1(_03871_),
    .Y(_04034_));
 sky130_fd_sc_hd__or3_1 _09642_ (.A(_04024_),
    .B(_04030_),
    .C(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__o21ai_1 _09643_ (.A1(_04030_),
    .A2(_04034_),
    .B1(_04024_),
    .Y(_04036_));
 sky130_fd_sc_hd__nand2_1 _09644_ (.A(_04035_),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__or3b_1 _09645_ (.A(_03998_),
    .B(_04022_),
    .C_N(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__o21bai_1 _09646_ (.A1(_03998_),
    .A2(_04022_),
    .B1_N(_04037_),
    .Y(_04039_));
 sky130_fd_sc_hd__or2b_1 _09647_ (.A(_04015_),
    .B_N(_04017_),
    .X(_04040_));
 sky130_fd_sc_hd__o21ai_1 _09648_ (.A1(_03996_),
    .A2(_04018_),
    .B1(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__and3_1 _09649_ (.A(_04038_),
    .B(_04039_),
    .C(_04041_),
    .X(_04042_));
 sky130_fd_sc_hd__a21oi_1 _09650_ (.A1(_04038_),
    .A2(_04039_),
    .B1(_04041_),
    .Y(_04043_));
 sky130_fd_sc_hd__o21ai_1 _09651_ (.A1(_04042_),
    .A2(_04043_),
    .B1(_03868_),
    .Y(_04044_));
 sky130_fd_sc_hd__o211a_1 _09652_ (.A1(\_185_[5] ),
    .A2(_03869_),
    .B1(_03919_),
    .C1(_04044_),
    .X(_00414_));
 sky130_fd_sc_hd__or2_1 _09653_ (.A(\_243_[6] ),
    .B(_03914_),
    .X(_04045_));
 sky130_fd_sc_hd__o22a_1 _09654_ (.A1(\_246_[6] ),
    .A2(_01313_),
    .B1(_01299_),
    .B2(\_179_[6] ),
    .X(_04046_));
 sky130_fd_sc_hd__and3_1 _09655_ (.A(\_142_[6] ),
    .B(_04045_),
    .C(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__a21oi_1 _09656_ (.A1(_04045_),
    .A2(_04046_),
    .B1(\_142_[6] ),
    .Y(_04048_));
 sky130_fd_sc_hd__or2_1 _09657_ (.A(_04047_),
    .B(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__nand2_1 _09658_ (.A(_03957_),
    .B(_03887_),
    .Y(_04050_));
 sky130_fd_sc_hd__nand2_2 _09659_ (.A(_01278_),
    .B(_01292_),
    .Y(_04051_));
 sky130_fd_sc_hd__a31o_1 _09660_ (.A1(_03884_),
    .A2(_04051_),
    .A3(_03925_),
    .B1(_03930_),
    .X(_04052_));
 sky130_fd_sc_hd__a21bo_1 _09661_ (.A1(_04028_),
    .A2(_04050_),
    .B1_N(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__nor2_1 _09662_ (.A(_01230_),
    .B(_03933_),
    .Y(_04054_));
 sky130_fd_sc_hd__nor2_2 _09663_ (.A(_01241_),
    .B(_01280_),
    .Y(_04055_));
 sky130_fd_sc_hd__nand2_1 _09664_ (.A(_01284_),
    .B(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__nand2_1 _09665_ (.A(_03884_),
    .B(_03901_),
    .Y(_04057_));
 sky130_fd_sc_hd__and3_1 _09666_ (.A(_03890_),
    .B(_03896_),
    .C(_03898_),
    .X(_04058_));
 sky130_fd_sc_hd__or2_1 _09667_ (.A(_03884_),
    .B(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__nor2_2 _09668_ (.A(_01230_),
    .B(_01235_),
    .Y(_04060_));
 sky130_fd_sc_hd__o211a_1 _09669_ (.A1(_01292_),
    .A2(_04057_),
    .B1(_04059_),
    .C1(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__a221o_1 _09670_ (.A1(_03871_),
    .A2(_04053_),
    .B1(_04054_),
    .B2(_04056_),
    .C1(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__xor2_1 _09671_ (.A(_04049_),
    .B(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__a21bo_1 _09672_ (.A1(\_142_[5] ),
    .A2(_04023_),
    .B1_N(_04035_),
    .X(_04064_));
 sky130_fd_sc_hd__xnor2_1 _09673_ (.A(_04063_),
    .B(_04064_),
    .Y(_04065_));
 sky130_fd_sc_hd__inv_2 _09674_ (.A(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__inv_2 _09675_ (.A(_04038_),
    .Y(_04067_));
 sky130_fd_sc_hd__o211a_1 _09676_ (.A1(_03996_),
    .A2(_04018_),
    .B1(_04039_),
    .C1(_04040_),
    .X(_04068_));
 sky130_fd_sc_hd__or2_1 _09677_ (.A(_04067_),
    .B(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__xnor2_1 _09678_ (.A(_04066_),
    .B(_04069_),
    .Y(_04070_));
 sky130_fd_sc_hd__nand2_1 _09679_ (.A(_03870_),
    .B(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__o211a_1 _09680_ (.A1(\_185_[6] ),
    .A2(_03869_),
    .B1(_03919_),
    .C1(_04071_),
    .X(_00415_));
 sky130_fd_sc_hd__and2b_1 _09681_ (.A_N(_04049_),
    .B(_04062_),
    .X(_04072_));
 sky130_fd_sc_hd__o221a_1 _09682_ (.A1(\_246_[7] ),
    .A2(_01314_),
    .B1(_03914_),
    .B2(\_243_[7] ),
    .C1(_01452_),
    .X(_04073_));
 sky130_fd_sc_hd__xnor2_1 _09683_ (.A(\_142_[7] ),
    .B(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__buf_2 _09684_ (.A(_04002_),
    .X(_04075_));
 sky130_fd_sc_hd__or2_1 _09685_ (.A(_04002_),
    .B(_01278_),
    .X(_04076_));
 sky130_fd_sc_hd__nor2_1 _09686_ (.A(_03923_),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__clkbuf_4 _09687_ (.A(_03933_),
    .X(_04078_));
 sky130_fd_sc_hd__a311o_1 _09688_ (.A1(_04075_),
    .A2(_03954_),
    .A3(_03928_),
    .B1(_04077_),
    .C1(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__nand2_2 _09689_ (.A(_03896_),
    .B(_03888_),
    .Y(_04080_));
 sky130_fd_sc_hd__nand2_1 _09690_ (.A(_03884_),
    .B(_03898_),
    .Y(_04081_));
 sky130_fd_sc_hd__nor2_1 _09691_ (.A(_01278_),
    .B(_03878_),
    .Y(_04082_));
 sky130_fd_sc_hd__nor2_1 _09692_ (.A(_04081_),
    .B(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__a211o_1 _09693_ (.A1(_04075_),
    .A2(_04080_),
    .B1(_04083_),
    .C1(_03872_),
    .X(_04084_));
 sky130_fd_sc_hd__nand2_1 _09694_ (.A(_03884_),
    .B(_03927_),
    .Y(_04085_));
 sky130_fd_sc_hd__or4_1 _09695_ (.A(_01235_),
    .B(_03875_),
    .C(_04005_),
    .D(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__nor2_2 _09696_ (.A(_01241_),
    .B(_01283_),
    .Y(_04087_));
 sky130_fd_sc_hd__and4_1 _09697_ (.A(_01234_),
    .B(_03884_),
    .C(_03903_),
    .D(_03928_),
    .X(_04088_));
 sky130_fd_sc_hd__a21oi_1 _09698_ (.A1(_03983_),
    .A2(_04087_),
    .B1(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__a21oi_1 _09699_ (.A1(_04086_),
    .A2(_04089_),
    .B1(_03871_),
    .Y(_04090_));
 sky130_fd_sc_hd__a31o_1 _09700_ (.A1(_01231_),
    .A2(_04079_),
    .A3(_04084_),
    .B1(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__xor2_1 _09701_ (.A(_04074_),
    .B(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__o21ai_1 _09702_ (.A1(_04047_),
    .A2(_04072_),
    .B1(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__or3_1 _09703_ (.A(_04047_),
    .B(_04072_),
    .C(_04092_),
    .X(_04094_));
 sky130_fd_sc_hd__nand2_1 _09704_ (.A(_04093_),
    .B(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__or2b_1 _09705_ (.A(_04063_),
    .B_N(_04064_),
    .X(_04096_));
 sky130_fd_sc_hd__o21ai_1 _09706_ (.A1(_04066_),
    .A2(_04069_),
    .B1(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__o21ai_1 _09707_ (.A1(_04095_),
    .A2(_04097_),
    .B1(_03867_),
    .Y(_04098_));
 sky130_fd_sc_hd__a21o_1 _09708_ (.A1(_04095_),
    .A2(_04097_),
    .B1(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__o211a_1 _09709_ (.A1(\_185_[7] ),
    .A2(_03869_),
    .B1(_03919_),
    .C1(_04099_),
    .X(_00416_));
 sky130_fd_sc_hd__nor2_1 _09710_ (.A(_04074_),
    .B(_04091_),
    .Y(_04100_));
 sky130_fd_sc_hd__a21oi_1 _09711_ (.A1(\_142_[7] ),
    .A2(_04073_),
    .B1(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__or2_1 _09712_ (.A(_03886_),
    .B(_04025_),
    .X(_04102_));
 sky130_fd_sc_hd__nand2_2 _09713_ (.A(_04002_),
    .B(_03901_),
    .Y(_04103_));
 sky130_fd_sc_hd__or2_1 _09714_ (.A(_04103_),
    .B(_04080_),
    .X(_04104_));
 sky130_fd_sc_hd__a221oi_1 _09715_ (.A1(_01281_),
    .A2(_03960_),
    .B1(_04080_),
    .B2(_04075_),
    .C1(_03872_),
    .Y(_04105_));
 sky130_fd_sc_hd__a31o_1 _09716_ (.A1(_01236_),
    .A2(_04102_),
    .A3(_04104_),
    .B1(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__nand2_2 _09717_ (.A(_01242_),
    .B(_03890_),
    .Y(_04107_));
 sky130_fd_sc_hd__or2_1 _09718_ (.A(_04002_),
    .B(_01283_),
    .X(_04108_));
 sky130_fd_sc_hd__o2111a_1 _09719_ (.A1(_03886_),
    .A2(_04103_),
    .B1(_04107_),
    .C1(_04108_),
    .D1(_04054_),
    .X(_04109_));
 sky130_fd_sc_hd__or2_1 _09720_ (.A(_04081_),
    .B(_04010_),
    .X(_04110_));
 sky130_fd_sc_hd__o311a_1 _09721_ (.A1(_01242_),
    .A2(_03897_),
    .A3(_04031_),
    .B1(_04110_),
    .C1(_04060_),
    .X(_04111_));
 sky130_fd_sc_hd__a211o_1 _09722_ (.A1(_01231_),
    .A2(_04106_),
    .B1(_04109_),
    .C1(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__o221a_1 _09723_ (.A1(\_246_[8] ),
    .A2(_01314_),
    .B1(_03914_),
    .B2(\_243_[8] ),
    .C1(_01455_),
    .X(_04113_));
 sky130_fd_sc_hd__and2_1 _09724_ (.A(\_142_[8] ),
    .B(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__nor2_1 _09725_ (.A(\_142_[8] ),
    .B(_04113_),
    .Y(_04115_));
 sky130_fd_sc_hd__or2_1 _09726_ (.A(_04114_),
    .B(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__nor2_1 _09727_ (.A(_04112_),
    .B(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__and2_1 _09728_ (.A(_04112_),
    .B(_04116_),
    .X(_04118_));
 sky130_fd_sc_hd__nor2_1 _09729_ (.A(_04117_),
    .B(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__and2b_1 _09730_ (.A_N(_04101_),
    .B(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__and2b_1 _09731_ (.A_N(_04119_),
    .B(_04101_),
    .X(_04121_));
 sky130_fd_sc_hd__or2_1 _09732_ (.A(_04120_),
    .B(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__a21bo_1 _09733_ (.A1(_04096_),
    .A2(_04093_),
    .B1_N(_04094_),
    .X(_04123_));
 sky130_fd_sc_hd__o41ai_2 _09734_ (.A1(_04067_),
    .A2(_04066_),
    .A3(_04068_),
    .A4(_04095_),
    .B1(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__and2b_1 _09735_ (.A_N(_04122_),
    .B(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__and2b_1 _09736_ (.A_N(_04124_),
    .B(_04122_),
    .X(_04126_));
 sky130_fd_sc_hd__o21ai_1 _09737_ (.A1(_04125_),
    .A2(_04126_),
    .B1(_03868_),
    .Y(_04127_));
 sky130_fd_sc_hd__o211a_1 _09738_ (.A1(\_185_[8] ),
    .A2(_03869_),
    .B1(_03919_),
    .C1(_04127_),
    .X(_00417_));
 sky130_fd_sc_hd__nor2_1 _09739_ (.A(_04120_),
    .B(_04125_),
    .Y(_04128_));
 sky130_fd_sc_hd__buf_2 _09740_ (.A(_03914_),
    .X(_04129_));
 sky130_fd_sc_hd__o221a_1 _09741_ (.A1(\_246_[9] ),
    .A2(_01314_),
    .B1(_04129_),
    .B2(\_243_[9] ),
    .C1(_01457_),
    .X(_04130_));
 sky130_fd_sc_hd__xnor2_1 _09742_ (.A(\_142_[9] ),
    .B(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__clkbuf_4 _09743_ (.A(_03961_),
    .X(_04132_));
 sky130_fd_sc_hd__or3_1 _09744_ (.A(_03933_),
    .B(_04087_),
    .C(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__or3_1 _09745_ (.A(_03886_),
    .B(_04010_),
    .C(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__a31oi_1 _09746_ (.A1(_01242_),
    .A2(_03890_),
    .A3(_03898_),
    .B1(_03872_),
    .Y(_04135_));
 sky130_fd_sc_hd__a21oi_1 _09747_ (.A1(_04056_),
    .A2(_04135_),
    .B1(_01231_),
    .Y(_04136_));
 sky130_fd_sc_hd__o211a_1 _09748_ (.A1(_04080_),
    .A2(_04107_),
    .B1(_04050_),
    .C1(_03872_),
    .X(_04137_));
 sky130_fd_sc_hd__nor2_1 _09749_ (.A(_01284_),
    .B(_03903_),
    .Y(_04138_));
 sky130_fd_sc_hd__nand2_1 _09750_ (.A(_01242_),
    .B(_03873_),
    .Y(_04139_));
 sky130_fd_sc_hd__o221a_1 _09751_ (.A1(_04103_),
    .A2(_04010_),
    .B1(_04138_),
    .B2(_04139_),
    .C1(_04078_),
    .X(_04140_));
 sky130_fd_sc_hd__nor2_1 _09752_ (.A(_04137_),
    .B(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__a22o_1 _09753_ (.A1(_04134_),
    .A2(_04136_),
    .B1(_04141_),
    .B2(_01231_),
    .X(_04142_));
 sky130_fd_sc_hd__xor2_1 _09754_ (.A(_04131_),
    .B(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__or3_1 _09755_ (.A(_04114_),
    .B(_04117_),
    .C(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__o21a_1 _09756_ (.A1(_04114_),
    .A2(_04117_),
    .B1(_04143_),
    .X(_04145_));
 sky130_fd_sc_hd__inv_2 _09757_ (.A(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__nand2_1 _09758_ (.A(_04144_),
    .B(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__xnor2_1 _09759_ (.A(_04128_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__nand2_1 _09760_ (.A(_03868_),
    .B(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__o211a_1 _09761_ (.A1(\_185_[9] ),
    .A2(_03869_),
    .B1(_03919_),
    .C1(_04149_),
    .X(_00418_));
 sky130_fd_sc_hd__buf_2 _09762_ (.A(_03868_),
    .X(_04150_));
 sky130_fd_sc_hd__nand2_1 _09763_ (.A(_04128_),
    .B(_04146_),
    .Y(_04151_));
 sky130_fd_sc_hd__o221a_1 _09764_ (.A1(\_246_[10] ),
    .A2(_01314_),
    .B1(_03914_),
    .B2(\_243_[10] ),
    .C1(_01462_),
    .X(_04152_));
 sky130_fd_sc_hd__and2_1 _09765_ (.A(\_142_[10] ),
    .B(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__nor2_1 _09766_ (.A(\_142_[10] ),
    .B(_04152_),
    .Y(_04154_));
 sky130_fd_sc_hd__or2_1 _09767_ (.A(_04153_),
    .B(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__nor2_1 _09768_ (.A(_01243_),
    .B(_03983_),
    .Y(_04156_));
 sky130_fd_sc_hd__nand2_1 _09769_ (.A(_03910_),
    .B(_01236_),
    .Y(_04157_));
 sky130_fd_sc_hd__nor2_1 _09770_ (.A(_03934_),
    .B(_04005_),
    .Y(_04158_));
 sky130_fd_sc_hd__a211o_1 _09771_ (.A1(_04156_),
    .A2(_03925_),
    .B1(_04157_),
    .C1(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__nor2_1 _09772_ (.A(_04075_),
    .B(_03897_),
    .Y(_04160_));
 sky130_fd_sc_hd__or2_1 _09773_ (.A(_01230_),
    .B(_03872_),
    .X(_04161_));
 sky130_fd_sc_hd__a221o_1 _09774_ (.A1(_04051_),
    .A2(_04132_),
    .B1(_04160_),
    .B2(_03903_),
    .C1(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__o21a_1 _09775_ (.A1(_04010_),
    .A2(_03936_),
    .B1(_04002_),
    .X(_04163_));
 sky130_fd_sc_hd__nand2_1 _09776_ (.A(_03872_),
    .B(_04057_),
    .Y(_04164_));
 sky130_fd_sc_hd__a32o_1 _09777_ (.A1(_03884_),
    .A2(_03898_),
    .A3(_03873_),
    .B1(_04006_),
    .B2(_04051_),
    .X(_04165_));
 sky130_fd_sc_hd__o22a_1 _09778_ (.A1(_04163_),
    .A2(_04164_),
    .B1(_04165_),
    .B2(_03872_),
    .X(_04166_));
 sky130_fd_sc_hd__or2_1 _09779_ (.A(_03910_),
    .B(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__and3_1 _09780_ (.A(_04159_),
    .B(_04162_),
    .C(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__xnor2_1 _09781_ (.A(_04155_),
    .B(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__o2bb2ai_1 _09782_ (.A1_N(\_142_[9] ),
    .A2_N(_04130_),
    .B1(_04131_),
    .B2(_04142_),
    .Y(_04170_));
 sky130_fd_sc_hd__xnor2_1 _09783_ (.A(_04169_),
    .B(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__a21oi_1 _09784_ (.A1(_04144_),
    .A2(_04151_),
    .B1(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__and3_1 _09785_ (.A(_04144_),
    .B(_04151_),
    .C(_04171_),
    .X(_04173_));
 sky130_fd_sc_hd__o21ai_1 _09786_ (.A1(_04172_),
    .A2(_04173_),
    .B1(_03868_),
    .Y(_04174_));
 sky130_fd_sc_hd__o211a_1 _09787_ (.A1(\_185_[10] ),
    .A2(_04150_),
    .B1(_03919_),
    .C1(_04174_),
    .X(_00419_));
 sky130_fd_sc_hd__buf_2 _09788_ (.A(_02833_),
    .X(_04175_));
 sky130_fd_sc_hd__nor2_1 _09789_ (.A(_04155_),
    .B(_04168_),
    .Y(_04176_));
 sky130_fd_sc_hd__nand2_1 _09790_ (.A(_01283_),
    .B(_03952_),
    .Y(_04177_));
 sky130_fd_sc_hd__o311a_1 _09791_ (.A1(_04002_),
    .A2(_01292_),
    .A3(_04027_),
    .B1(_04177_),
    .C1(_01235_),
    .X(_04178_));
 sky130_fd_sc_hd__nor2_1 _09792_ (.A(_03934_),
    .B(_03923_),
    .Y(_04179_));
 sky130_fd_sc_hd__a211oi_1 _09793_ (.A1(_03954_),
    .A2(_03876_),
    .B1(_04179_),
    .C1(_01235_),
    .Y(_04180_));
 sky130_fd_sc_hd__a21oi_1 _09794_ (.A1(_03898_),
    .A2(_03893_),
    .B1(_03876_),
    .Y(_04181_));
 sky130_fd_sc_hd__nor2_1 _09795_ (.A(_03933_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__a22o_1 _09796_ (.A1(_04055_),
    .A2(_04080_),
    .B1(_03928_),
    .B2(_03880_),
    .X(_04183_));
 sky130_fd_sc_hd__o21ai_1 _09797_ (.A1(_03872_),
    .A2(_04183_),
    .B1(_01230_),
    .Y(_04184_));
 sky130_fd_sc_hd__o32a_1 _09798_ (.A1(_01230_),
    .A2(_04178_),
    .A3(_04180_),
    .B1(_04182_),
    .B2(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__inv_2 _09799_ (.A(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__o221a_1 _09800_ (.A1(\_246_[11] ),
    .A2(_01314_),
    .B1(_03914_),
    .B2(\_243_[11] ),
    .C1(_01464_),
    .X(_04187_));
 sky130_fd_sc_hd__and2_1 _09801_ (.A(\_142_[11] ),
    .B(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__nor2_1 _09802_ (.A(\_142_[11] ),
    .B(_04187_),
    .Y(_04189_));
 sky130_fd_sc_hd__or2_1 _09803_ (.A(_04188_),
    .B(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__nor2_1 _09804_ (.A(_04186_),
    .B(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__and2_1 _09805_ (.A(_04186_),
    .B(_04190_),
    .X(_04192_));
 sky130_fd_sc_hd__or2_1 _09806_ (.A(_04191_),
    .B(_04192_),
    .X(_04193_));
 sky130_fd_sc_hd__or3b_1 _09807_ (.A(_04153_),
    .B(_04176_),
    .C_N(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__o21bai_2 _09808_ (.A1(_04153_),
    .A2(_04176_),
    .B1_N(_04193_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_1 _09809_ (.A(_04194_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__and2b_1 _09810_ (.A_N(_04169_),
    .B(_04170_),
    .X(_04197_));
 sky130_fd_sc_hd__a31o_1 _09811_ (.A1(_04144_),
    .A2(_04151_),
    .A3(_04171_),
    .B1(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__xor2_1 _09812_ (.A(_04196_),
    .B(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__nand2_1 _09813_ (.A(_03868_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__o211a_1 _09814_ (.A1(\_185_[11] ),
    .A2(_04150_),
    .B1(_04175_),
    .C1(_04200_),
    .X(_00420_));
 sky130_fd_sc_hd__nand3_1 _09815_ (.A(_04171_),
    .B(_04194_),
    .C(_04195_),
    .Y(_04201_));
 sky130_fd_sc_hd__or4b_1 _09816_ (.A(_04122_),
    .B(_04147_),
    .C(_04201_),
    .D_N(_04124_),
    .X(_04202_));
 sky130_fd_sc_hd__o21ai_1 _09817_ (.A1(_04120_),
    .A2(_04145_),
    .B1(_04144_),
    .Y(_04203_));
 sky130_fd_sc_hd__o2bb2a_1 _09818_ (.A1_N(_04197_),
    .A2_N(_04194_),
    .B1(_04201_),
    .B2(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__and3_1 _09819_ (.A(_04195_),
    .B(_04202_),
    .C(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__o221a_1 _09820_ (.A1(\_246_[12] ),
    .A2(_01314_),
    .B1(_03914_),
    .B2(\_243_[12] ),
    .C1(_01466_),
    .X(_04206_));
 sky130_fd_sc_hd__and2_1 _09821_ (.A(\_142_[12] ),
    .B(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__nor2_1 _09822_ (.A(\_142_[12] ),
    .B(_04206_),
    .Y(_04208_));
 sky130_fd_sc_hd__nor2_1 _09823_ (.A(_04207_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__clkbuf_4 _09824_ (.A(_03910_),
    .X(_04210_));
 sky130_fd_sc_hd__a311o_1 _09825_ (.A1(_01242_),
    .A2(_03883_),
    .A3(_03984_),
    .B1(_04055_),
    .C1(_03876_),
    .X(_04211_));
 sky130_fd_sc_hd__nand2_1 _09826_ (.A(_01236_),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__a221o_1 _09827_ (.A1(_03898_),
    .A2(_03880_),
    .B1(_04132_),
    .B2(_03888_),
    .C1(_01236_),
    .X(_04213_));
 sky130_fd_sc_hd__a32o_1 _09828_ (.A1(_01242_),
    .A2(_01280_),
    .A3(_04080_),
    .B1(_04087_),
    .B2(_03983_),
    .X(_04214_));
 sky130_fd_sc_hd__a21o_1 _09829_ (.A1(_04002_),
    .A2(_04005_),
    .B1(_03933_),
    .X(_04215_));
 sky130_fd_sc_hd__a41o_1 _09830_ (.A1(_01242_),
    .A2(_03890_),
    .A3(_03896_),
    .A4(_03927_),
    .B1(_04215_),
    .X(_04216_));
 sky130_fd_sc_hd__o211a_1 _09831_ (.A1(_01236_),
    .A2(_04214_),
    .B1(_04216_),
    .C1(_03871_),
    .X(_04217_));
 sky130_fd_sc_hd__a31o_1 _09832_ (.A1(_04210_),
    .A2(_04212_),
    .A3(_04213_),
    .B1(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__and2_1 _09833_ (.A(_04209_),
    .B(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__nor2_1 _09834_ (.A(_04209_),
    .B(_04218_),
    .Y(_04220_));
 sky130_fd_sc_hd__or2_1 _09835_ (.A(_04219_),
    .B(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__o21bai_2 _09836_ (.A1(_04188_),
    .A2(_04191_),
    .B1_N(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__or3b_1 _09837_ (.A(_04188_),
    .B(_04191_),
    .C_N(_04221_),
    .X(_04223_));
 sky130_fd_sc_hd__nand2_1 _09838_ (.A(_04222_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__or2_1 _09839_ (.A(_04205_),
    .B(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__nand2_1 _09840_ (.A(_04205_),
    .B(_04224_),
    .Y(_04226_));
 sky130_fd_sc_hd__a21o_1 _09841_ (.A1(_04225_),
    .A2(_04226_),
    .B1(_03946_),
    .X(_04227_));
 sky130_fd_sc_hd__o211a_1 _09842_ (.A1(\_185_[12] ),
    .A2(_04150_),
    .B1(_04175_),
    .C1(_04227_),
    .X(_00421_));
 sky130_fd_sc_hd__o221a_1 _09843_ (.A1(\_246_[13] ),
    .A2(_01315_),
    .B1(_04129_),
    .B2(\_243_[13] ),
    .C1(_01469_),
    .X(_04228_));
 sky130_fd_sc_hd__xnor2_1 _09844_ (.A(\_142_[13] ),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand2_1 _09845_ (.A(_03896_),
    .B(_03927_),
    .Y(_04230_));
 sky130_fd_sc_hd__or2_1 _09846_ (.A(_01242_),
    .B(_04230_),
    .X(_04231_));
 sky130_fd_sc_hd__a211oi_1 _09847_ (.A1(_01281_),
    .A2(_04231_),
    .B1(_03908_),
    .C1(_01231_),
    .Y(_04232_));
 sky130_fd_sc_hd__or2_1 _09848_ (.A(_04087_),
    .B(_03958_),
    .X(_04233_));
 sky130_fd_sc_hd__a31o_1 _09849_ (.A1(_03871_),
    .A2(_03925_),
    .A3(_04233_),
    .B1(_04078_),
    .X(_04234_));
 sky130_fd_sc_hd__and2_1 _09850_ (.A(_03905_),
    .B(_03981_),
    .X(_04235_));
 sky130_fd_sc_hd__o21a_1 _09851_ (.A1(_01283_),
    .A2(_03958_),
    .B1(_03904_),
    .X(_04236_));
 sky130_fd_sc_hd__or3_1 _09852_ (.A(_03910_),
    .B(_03906_),
    .C(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__o31a_1 _09853_ (.A1(_03871_),
    .A2(_03897_),
    .A3(_04235_),
    .B1(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__o22a_1 _09854_ (.A1(_04232_),
    .A2(_04234_),
    .B1(_04238_),
    .B2(_01237_),
    .X(_04239_));
 sky130_fd_sc_hd__nor2_1 _09855_ (.A(_04229_),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__and2_1 _09856_ (.A(_04229_),
    .B(_04239_),
    .X(_04241_));
 sky130_fd_sc_hd__or2_1 _09857_ (.A(_04240_),
    .B(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__o21ba_1 _09858_ (.A1(_04207_),
    .A2(_04219_),
    .B1_N(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__or3b_1 _09859_ (.A(_04207_),
    .B(_04219_),
    .C_N(_04242_),
    .X(_04244_));
 sky130_fd_sc_hd__and2b_1 _09860_ (.A_N(_04243_),
    .B(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__and3_1 _09861_ (.A(_04222_),
    .B(_04225_),
    .C(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__a21oi_1 _09862_ (.A1(_04222_),
    .A2(_04225_),
    .B1(_04245_),
    .Y(_04247_));
 sky130_fd_sc_hd__or3_1 _09863_ (.A(_03945_),
    .B(_04246_),
    .C(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__o211a_1 _09864_ (.A1(\_185_[13] ),
    .A2(_04150_),
    .B1(_04175_),
    .C1(_04248_),
    .X(_00422_));
 sky130_fd_sc_hd__o221a_1 _09865_ (.A1(\_246_[14] ),
    .A2(_01314_),
    .B1(_04129_),
    .B2(\_243_[14] ),
    .C1(_01472_),
    .X(_04249_));
 sky130_fd_sc_hd__and2_1 _09866_ (.A(\_142_[14] ),
    .B(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__nor2_1 _09867_ (.A(\_142_[14] ),
    .B(_04249_),
    .Y(_04251_));
 sky130_fd_sc_hd__nor2_1 _09868_ (.A(_04250_),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand2_1 _09869_ (.A(_03880_),
    .B(_03927_),
    .Y(_04253_));
 sky130_fd_sc_hd__o31a_1 _09870_ (.A1(_01243_),
    .A2(_04010_),
    .A3(_03936_),
    .B1(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__nand2_1 _09871_ (.A(_01231_),
    .B(_01236_),
    .Y(_04255_));
 sky130_fd_sc_hd__a21o_1 _09872_ (.A1(_04103_),
    .A2(_04110_),
    .B1(_03935_),
    .X(_04256_));
 sky130_fd_sc_hd__or4_1 _09873_ (.A(_03871_),
    .B(_04078_),
    .C(_04132_),
    .D(_04058_),
    .X(_04257_));
 sky130_fd_sc_hd__and3_1 _09874_ (.A(_04002_),
    .B(_03888_),
    .C(_03929_),
    .X(_04258_));
 sky130_fd_sc_hd__or4_1 _09875_ (.A(_03910_),
    .B(_01236_),
    .C(_04179_),
    .D(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__o211a_1 _09876_ (.A1(_04255_),
    .A2(_04256_),
    .B1(_04257_),
    .C1(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__o21ai_1 _09877_ (.A1(_04161_),
    .A2(_04254_),
    .B1(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__and2_1 _09878_ (.A(_04252_),
    .B(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__nor2_1 _09879_ (.A(_04252_),
    .B(_04261_),
    .Y(_04263_));
 sky130_fd_sc_hd__or2_1 _09880_ (.A(_04262_),
    .B(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__a21oi_1 _09881_ (.A1(\_142_[13] ),
    .A2(_04228_),
    .B1(_04240_),
    .Y(_04265_));
 sky130_fd_sc_hd__xnor2_1 _09882_ (.A(_04264_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__or3b_1 _09883_ (.A(_04224_),
    .B(_04243_),
    .C_N(_04244_),
    .X(_04267_));
 sky130_fd_sc_hd__inv_2 _09884_ (.A(_04222_),
    .Y(_04268_));
 sky130_fd_sc_hd__o21ai_1 _09885_ (.A1(_04268_),
    .A2(_04243_),
    .B1(_04244_),
    .Y(_04269_));
 sky130_fd_sc_hd__o21a_1 _09886_ (.A1(_04205_),
    .A2(_04267_),
    .B1(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__nand2_1 _09887_ (.A(_04266_),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__or2_1 _09888_ (.A(_04266_),
    .B(_04270_),
    .X(_04272_));
 sky130_fd_sc_hd__a21o_1 _09889_ (.A1(_04271_),
    .A2(_04272_),
    .B1(_03946_),
    .X(_04273_));
 sky130_fd_sc_hd__o211a_1 _09890_ (.A1(\_185_[14] ),
    .A2(_04150_),
    .B1(_04175_),
    .C1(_04273_),
    .X(_00423_));
 sky130_fd_sc_hd__o221a_1 _09891_ (.A1(\_246_[15] ),
    .A2(_01314_),
    .B1(_04129_),
    .B2(\_243_[15] ),
    .C1(_01475_),
    .X(_04274_));
 sky130_fd_sc_hd__and2_1 _09892_ (.A(\_142_[15] ),
    .B(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__nor2_1 _09893_ (.A(\_142_[15] ),
    .B(_04274_),
    .Y(_04276_));
 sky130_fd_sc_hd__or2_1 _09894_ (.A(_04275_),
    .B(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__o31a_1 _09895_ (.A1(_01242_),
    .A2(_04082_),
    .A3(_03936_),
    .B1(_01236_),
    .X(_04278_));
 sky130_fd_sc_hd__or2b_1 _09896_ (.A(_04011_),
    .B_N(_04278_),
    .X(_04279_));
 sky130_fd_sc_hd__nand2_1 _09897_ (.A(_04078_),
    .B(_04231_),
    .Y(_04280_));
 sky130_fd_sc_hd__a21o_1 _09898_ (.A1(_03905_),
    .A2(_04230_),
    .B1(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__a221o_1 _09899_ (.A1(_03888_),
    .A2(_04006_),
    .B1(_04080_),
    .B2(_01243_),
    .C1(_01237_),
    .X(_04282_));
 sky130_fd_sc_hd__o211a_1 _09900_ (.A1(_03886_),
    .A2(_03907_),
    .B1(_04139_),
    .C1(_01237_),
    .X(_04283_));
 sky130_fd_sc_hd__nor2_1 _09901_ (.A(_01231_),
    .B(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__a32o_1 _09902_ (.A1(_01232_),
    .A2(_04279_),
    .A3(_04281_),
    .B1(_04282_),
    .B2(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__xor2_1 _09903_ (.A(_04277_),
    .B(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__nor3_1 _09904_ (.A(_04250_),
    .B(_04262_),
    .C(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__o21ai_1 _09905_ (.A1(_04250_),
    .A2(_04262_),
    .B1(_04286_),
    .Y(_04288_));
 sky130_fd_sc_hd__or2b_1 _09906_ (.A(_04287_),
    .B_N(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__or2_1 _09907_ (.A(_04264_),
    .B(_04265_),
    .X(_04290_));
 sky130_fd_sc_hd__o21ai_1 _09908_ (.A1(_04266_),
    .A2(_04270_),
    .B1(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__a21oi_1 _09909_ (.A1(_04289_),
    .A2(_04291_),
    .B1(_03945_),
    .Y(_04292_));
 sky130_fd_sc_hd__o21ai_1 _09910_ (.A1(_04289_),
    .A2(_04291_),
    .B1(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__o211a_1 _09911_ (.A1(\_185_[15] ),
    .A2(_04150_),
    .B1(_04175_),
    .C1(_04293_),
    .X(_00424_));
 sky130_fd_sc_hd__or2_1 _09912_ (.A(_04266_),
    .B(_04289_),
    .X(_04294_));
 sky130_fd_sc_hd__o221a_1 _09913_ (.A1(_04290_),
    .A2(_04287_),
    .B1(_04294_),
    .B2(_04269_),
    .C1(_04288_),
    .X(_04295_));
 sky130_fd_sc_hd__a311o_1 _09914_ (.A1(_04195_),
    .A2(_04202_),
    .A3(_04204_),
    .B1(_04267_),
    .C1(_04294_),
    .X(_04296_));
 sky130_fd_sc_hd__nor2_1 _09915_ (.A(_04277_),
    .B(_04285_),
    .Y(_04297_));
 sky130_fd_sc_hd__o221a_1 _09916_ (.A1(\_246_[16] ),
    .A2(_01315_),
    .B1(_04129_),
    .B2(\_243_[16] ),
    .C1(_01477_),
    .X(_04298_));
 sky130_fd_sc_hd__xnor2_1 _09917_ (.A(\_142_[16] ),
    .B(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__a211o_1 _09918_ (.A1(_03880_),
    .A2(_03984_),
    .B1(_04132_),
    .C1(_01237_),
    .X(_04300_));
 sky130_fd_sc_hd__o31a_1 _09919_ (.A1(_03983_),
    .A2(_04138_),
    .A3(_04133_),
    .B1(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__and2b_1 _09920_ (.A_N(_04011_),
    .B(_04231_),
    .X(_04302_));
 sky130_fd_sc_hd__nor2_2 _09921_ (.A(_01278_),
    .B(_01281_),
    .Y(_04303_));
 sky130_fd_sc_hd__or4_1 _09922_ (.A(_04075_),
    .B(_01285_),
    .C(_03875_),
    .D(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__or3b_1 _09923_ (.A(_01232_),
    .B(_04280_),
    .C_N(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__o221a_1 _09924_ (.A1(_04210_),
    .A2(_04301_),
    .B1(_04302_),
    .B2(_04157_),
    .C1(_04305_),
    .X(_04306_));
 sky130_fd_sc_hd__xnor2_1 _09925_ (.A(_04299_),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__o21bai_2 _09926_ (.A1(_04275_),
    .A2(_04297_),
    .B1_N(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__or3b_1 _09927_ (.A(_04275_),
    .B(_04297_),
    .C_N(_04307_),
    .X(_04309_));
 sky130_fd_sc_hd__nand2_1 _09928_ (.A(_04308_),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__a21o_1 _09929_ (.A1(_04295_),
    .A2(_04296_),
    .B1(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__nand3_1 _09930_ (.A(_04295_),
    .B(_04296_),
    .C(_04310_),
    .Y(_04312_));
 sky130_fd_sc_hd__a21o_1 _09931_ (.A1(_04311_),
    .A2(_04312_),
    .B1(_03945_),
    .X(_04313_));
 sky130_fd_sc_hd__o211a_1 _09932_ (.A1(\_185_[16] ),
    .A2(_04150_),
    .B1(_04175_),
    .C1(_04313_),
    .X(_00425_));
 sky130_fd_sc_hd__a32o_1 _09933_ (.A1(_01243_),
    .A2(_01281_),
    .A3(_03960_),
    .B1(_03888_),
    .B2(_04132_),
    .X(_04314_));
 sky130_fd_sc_hd__nor2_1 _09934_ (.A(_01237_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__nand2_1 _09935_ (.A(_04075_),
    .B(_03890_),
    .Y(_04316_));
 sky130_fd_sc_hd__a31o_1 _09936_ (.A1(_01237_),
    .A2(_04316_),
    .A3(_04253_),
    .B1(_01232_),
    .X(_04317_));
 sky130_fd_sc_hd__and3_1 _09937_ (.A(_01243_),
    .B(_01284_),
    .C(_03904_),
    .X(_04318_));
 sky130_fd_sc_hd__a21oi_1 _09938_ (.A1(_04075_),
    .A2(_04005_),
    .B1(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__nand2_1 _09939_ (.A(_01243_),
    .B(_03950_),
    .Y(_04320_));
 sky130_fd_sc_hd__nor2_1 _09940_ (.A(_01243_),
    .B(_03904_),
    .Y(_04321_));
 sky130_fd_sc_hd__a2bb2o_1 _09941_ (.A1_N(_03878_),
    .A2_N(_04320_),
    .B1(_01284_),
    .B2(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__mux2_1 _09942_ (.A0(_04319_),
    .A1(_04322_),
    .S(_01237_),
    .X(_04323_));
 sky130_fd_sc_hd__o22a_1 _09943_ (.A1(_04315_),
    .A2(_04317_),
    .B1(_04323_),
    .B2(_04210_),
    .X(_04324_));
 sky130_fd_sc_hd__o221a_1 _09944_ (.A1(\_246_[17] ),
    .A2(_01315_),
    .B1(_04129_),
    .B2(\_243_[17] ),
    .C1(_01482_),
    .X(_04325_));
 sky130_fd_sc_hd__xnor2_1 _09945_ (.A(\_142_[17] ),
    .B(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__xnor2_1 _09946_ (.A(_04324_),
    .B(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__a2bb2o_1 _09947_ (.A1_N(_04299_),
    .A2_N(_04306_),
    .B1(\_142_[16] ),
    .B2(_04298_),
    .X(_04328_));
 sky130_fd_sc_hd__xnor2_1 _09948_ (.A(_04327_),
    .B(_04328_),
    .Y(_04329_));
 sky130_fd_sc_hd__and3b_1 _09949_ (.A_N(_04329_),
    .B(_04311_),
    .C(_04308_),
    .X(_04330_));
 sky130_fd_sc_hd__a21boi_1 _09950_ (.A1(_04308_),
    .A2(_04311_),
    .B1_N(_04329_),
    .Y(_04331_));
 sky130_fd_sc_hd__or3_1 _09951_ (.A(_03945_),
    .B(_04330_),
    .C(_04331_),
    .X(_04332_));
 sky130_fd_sc_hd__o211a_1 _09952_ (.A1(\_185_[17] ),
    .A2(_04150_),
    .B1(_04175_),
    .C1(_04332_),
    .X(_00426_));
 sky130_fd_sc_hd__nor2_1 _09953_ (.A(_03960_),
    .B(_03907_),
    .Y(_04333_));
 sky130_fd_sc_hd__or3_1 _09954_ (.A(_04179_),
    .B(_04215_),
    .C(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__o311a_1 _09955_ (.A1(_01237_),
    .A2(_03876_),
    .A3(_04083_),
    .B1(_04334_),
    .C1(_01231_),
    .X(_04335_));
 sky130_fd_sc_hd__o311a_1 _09956_ (.A1(_01281_),
    .A2(_04087_),
    .A3(_04080_),
    .B1(_03938_),
    .C1(_04054_),
    .X(_04336_));
 sky130_fd_sc_hd__o311a_1 _09957_ (.A1(_01243_),
    .A2(_03897_),
    .A3(_04005_),
    .B1(_03925_),
    .C1(_04051_),
    .X(_04337_));
 sky130_fd_sc_hd__a211o_1 _09958_ (.A1(_01284_),
    .A2(_04321_),
    .B1(_04161_),
    .C1(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__or3b_2 _09959_ (.A(_04335_),
    .B(_04336_),
    .C_N(_04338_),
    .X(_04339_));
 sky130_fd_sc_hd__o221a_1 _09960_ (.A1(\_246_[18] ),
    .A2(_01315_),
    .B1(_04129_),
    .B2(\_243_[18] ),
    .C1(_01486_),
    .X(_04340_));
 sky130_fd_sc_hd__xnor2_1 _09961_ (.A(\_142_[18] ),
    .B(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__xor2_1 _09962_ (.A(_04339_),
    .B(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__inv_2 _09963_ (.A(_04326_),
    .Y(_04343_));
 sky130_fd_sc_hd__a22o_1 _09964_ (.A1(\_142_[17] ),
    .A2(_04325_),
    .B1(_04343_),
    .B2(_04324_),
    .X(_04344_));
 sky130_fd_sc_hd__nand2_1 _09965_ (.A(_04342_),
    .B(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__or2_1 _09966_ (.A(_04342_),
    .B(_04344_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _09967_ (.A(_04345_),
    .B(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hd__nand2_1 _09968_ (.A(_04327_),
    .B(_04328_),
    .Y(_04348_));
 sky130_fd_sc_hd__nor2_1 _09969_ (.A(_04327_),
    .B(_04328_),
    .Y(_04349_));
 sky130_fd_sc_hd__a31o_1 _09970_ (.A1(_04308_),
    .A2(_04311_),
    .A3(_04348_),
    .B1(_04349_),
    .X(_04350_));
 sky130_fd_sc_hd__nand2_1 _09971_ (.A(_04347_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__or2_1 _09972_ (.A(_04347_),
    .B(_04350_),
    .X(_04352_));
 sky130_fd_sc_hd__a21o_1 _09973_ (.A1(_04351_),
    .A2(_04352_),
    .B1(_03945_),
    .X(_04353_));
 sky130_fd_sc_hd__o211a_1 _09974_ (.A1(\_185_[18] ),
    .A2(_04150_),
    .B1(_04175_),
    .C1(_04353_),
    .X(_00427_));
 sky130_fd_sc_hd__or2_1 _09975_ (.A(\_243_[19] ),
    .B(_04129_),
    .X(_04354_));
 sky130_fd_sc_hd__o22a_1 _09976_ (.A1(\_246_[19] ),
    .A2(_01315_),
    .B1(_01300_),
    .B2(\_179_[19] ),
    .X(_04355_));
 sky130_fd_sc_hd__and3_1 _09977_ (.A(\_142_[19] ),
    .B(_04354_),
    .C(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__a21oi_1 _09978_ (.A1(_04354_),
    .A2(_04355_),
    .B1(\_142_[19] ),
    .Y(_04357_));
 sky130_fd_sc_hd__or2_1 _09979_ (.A(_04356_),
    .B(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__nor2_1 _09980_ (.A(_04082_),
    .B(_04320_),
    .Y(_04359_));
 sky130_fd_sc_hd__and2_1 _09981_ (.A(_03878_),
    .B(_04132_),
    .X(_04360_));
 sky130_fd_sc_hd__o21ai_1 _09982_ (.A1(_04075_),
    .A2(_03928_),
    .B1(_04078_),
    .Y(_04361_));
 sky130_fd_sc_hd__a31o_1 _09983_ (.A1(_03901_),
    .A2(_04006_),
    .A3(_03873_),
    .B1(_03910_),
    .X(_04362_));
 sky130_fd_sc_hd__nor2_1 _09984_ (.A(_04075_),
    .B(_01284_),
    .Y(_04363_));
 sky130_fd_sc_hd__a21oi_1 _09985_ (.A1(_03896_),
    .A2(_04132_),
    .B1(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__and2b_1 _09986_ (.A_N(_04010_),
    .B(_03952_),
    .X(_04365_));
 sky130_fd_sc_hd__nor2_1 _09987_ (.A(_01292_),
    .B(_04076_),
    .Y(_04366_));
 sky130_fd_sc_hd__or4_1 _09988_ (.A(_01231_),
    .B(_01236_),
    .C(_04365_),
    .D(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__o221a_1 _09989_ (.A1(_04361_),
    .A2(_04362_),
    .B1(_04364_),
    .B2(_04255_),
    .C1(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__o31a_1 _09990_ (.A1(_04157_),
    .A2(_04359_),
    .A3(_04360_),
    .B1(_04368_),
    .X(_04369_));
 sky130_fd_sc_hd__xnor2_1 _09991_ (.A(_04358_),
    .B(_04369_),
    .Y(_04370_));
 sky130_fd_sc_hd__o2bb2ai_1 _09992_ (.A1_N(\_142_[18] ),
    .A2_N(_04340_),
    .B1(_04341_),
    .B2(_04339_),
    .Y(_04371_));
 sky130_fd_sc_hd__xnor2_1 _09993_ (.A(_04370_),
    .B(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__and3_1 _09994_ (.A(_04345_),
    .B(_04352_),
    .C(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__a21oi_1 _09995_ (.A1(_04345_),
    .A2(_04352_),
    .B1(_04372_),
    .Y(_04374_));
 sky130_fd_sc_hd__or3_1 _09996_ (.A(_03945_),
    .B(_04373_),
    .C(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__o211a_1 _09997_ (.A1(\_185_[19] ),
    .A2(_04150_),
    .B1(_04175_),
    .C1(_04375_),
    .X(_00428_));
 sky130_fd_sc_hd__nor2_1 _09998_ (.A(_04358_),
    .B(_04369_),
    .Y(_04376_));
 sky130_fd_sc_hd__or2_1 _09999_ (.A(\_243_[20] ),
    .B(_04129_),
    .X(_04377_));
 sky130_fd_sc_hd__o22a_1 _10000_ (.A1(\_246_[20] ),
    .A2(_01315_),
    .B1(_01301_),
    .B2(\_179_[20] ),
    .X(_04378_));
 sky130_fd_sc_hd__and3_1 _10001_ (.A(\_142_[20] ),
    .B(_04377_),
    .C(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__a21oi_1 _10002_ (.A1(_04377_),
    .A2(_04378_),
    .B1(\_142_[20] ),
    .Y(_04380_));
 sky130_fd_sc_hd__or2_1 _10003_ (.A(_04379_),
    .B(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__nand2_1 _10004_ (.A(_04076_),
    .B(_04104_),
    .Y(_04382_));
 sky130_fd_sc_hd__nor2_1 _10005_ (.A(_01292_),
    .B(_04316_),
    .Y(_04383_));
 sky130_fd_sc_hd__a21o_1 _10006_ (.A1(_01244_),
    .A2(_01281_),
    .B1(_04383_),
    .X(_04384_));
 sky130_fd_sc_hd__nand2_1 _10007_ (.A(_03960_),
    .B(_03952_),
    .Y(_04385_));
 sky130_fd_sc_hd__nor2_1 _10008_ (.A(_04303_),
    .B(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__or2_1 _10009_ (.A(_03893_),
    .B(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__nor2_1 _10010_ (.A(_03876_),
    .B(_03893_),
    .Y(_04388_));
 sky130_fd_sc_hd__mux4_1 _10011_ (.A0(_04382_),
    .A1(_04384_),
    .A2(_04387_),
    .A3(_04388_),
    .S0(_04078_),
    .S1(_04210_),
    .X(_04389_));
 sky130_fd_sc_hd__nor2_1 _10012_ (.A(_04381_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__nand2_1 _10013_ (.A(_04381_),
    .B(_04389_),
    .Y(_04391_));
 sky130_fd_sc_hd__or2b_1 _10014_ (.A(_04390_),
    .B_N(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__o21ba_1 _10015_ (.A1(_04356_),
    .A2(_04376_),
    .B1_N(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__or3b_1 _10016_ (.A(_04356_),
    .B(_04376_),
    .C_N(_04392_),
    .X(_04394_));
 sky130_fd_sc_hd__or2b_1 _10017_ (.A(_04393_),
    .B_N(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__and3_1 _10018_ (.A(_04345_),
    .B(_04346_),
    .C(_04372_),
    .X(_04396_));
 sky130_fd_sc_hd__or3b_1 _10019_ (.A(_04310_),
    .B(_04329_),
    .C_N(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__a21o_1 _10020_ (.A1(_04295_),
    .A2(_04296_),
    .B1(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__inv_2 _10021_ (.A(_04345_),
    .Y(_04399_));
 sky130_fd_sc_hd__or2b_1 _10022_ (.A(_04371_),
    .B_N(_04370_),
    .X(_04400_));
 sky130_fd_sc_hd__a21oi_1 _10023_ (.A1(_04308_),
    .A2(_04348_),
    .B1(_04349_),
    .Y(_04401_));
 sky130_fd_sc_hd__and2b_1 _10024_ (.A_N(_04370_),
    .B(_04371_),
    .X(_04402_));
 sky130_fd_sc_hd__a221o_1 _10025_ (.A1(_04399_),
    .A2(_04400_),
    .B1(_04396_),
    .B2(_04401_),
    .C1(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__inv_2 _10026_ (.A(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__and2_1 _10027_ (.A(_04398_),
    .B(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__or2_1 _10028_ (.A(_04395_),
    .B(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__nand2_1 _10029_ (.A(_04395_),
    .B(_04405_),
    .Y(_04407_));
 sky130_fd_sc_hd__a21o_1 _10030_ (.A1(_04406_),
    .A2(_04407_),
    .B1(_03945_),
    .X(_04408_));
 sky130_fd_sc_hd__o211a_1 _10031_ (.A1(\_185_[20] ),
    .A2(_03870_),
    .B1(_04175_),
    .C1(_04408_),
    .X(_00429_));
 sky130_fd_sc_hd__buf_2 _10032_ (.A(_04129_),
    .X(_04409_));
 sky130_fd_sc_hd__o221a_1 _10033_ (.A1(\_246_[21] ),
    .A2(_01315_),
    .B1(_04409_),
    .B2(\_243_[21] ),
    .C1(_01493_),
    .X(_04410_));
 sky130_fd_sc_hd__and2_1 _10034_ (.A(\_142_[21] ),
    .B(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__nor2_1 _10035_ (.A(\_142_[21] ),
    .B(_04410_),
    .Y(_04412_));
 sky130_fd_sc_hd__or2_1 _10036_ (.A(_04411_),
    .B(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__a2111o_1 _10037_ (.A1(_01244_),
    .A2(_03878_),
    .B1(_03976_),
    .C1(_03897_),
    .D1(_01237_),
    .X(_04414_));
 sky130_fd_sc_hd__o31a_1 _10038_ (.A1(_04078_),
    .A2(_04032_),
    .A3(_04383_),
    .B1(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__and3_1 _10039_ (.A(_01244_),
    .B(_03928_),
    .C(_03929_),
    .X(_04416_));
 sky130_fd_sc_hd__or2_1 _10040_ (.A(_04280_),
    .B(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__or3b_1 _10041_ (.A(_01243_),
    .B(_01278_),
    .C_N(_03873_),
    .X(_04418_));
 sky130_fd_sc_hd__o311a_1 _10042_ (.A1(_03886_),
    .A2(_03983_),
    .A3(_04107_),
    .B1(_04418_),
    .C1(_01238_),
    .X(_04419_));
 sky130_fd_sc_hd__nor2_1 _10043_ (.A(_01232_),
    .B(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__a22o_1 _10044_ (.A1(_01232_),
    .A2(_04415_),
    .B1(_04417_),
    .B2(_04420_),
    .X(_04421_));
 sky130_fd_sc_hd__nor2_1 _10045_ (.A(_04413_),
    .B(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__and2_1 _10046_ (.A(_04413_),
    .B(_04421_),
    .X(_04423_));
 sky130_fd_sc_hd__nor2_1 _10047_ (.A(_04422_),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__o21a_1 _10048_ (.A1(_04379_),
    .A2(_04390_),
    .B1(_04424_),
    .X(_04425_));
 sky130_fd_sc_hd__or3_1 _10049_ (.A(_04379_),
    .B(_04390_),
    .C(_04424_),
    .X(_04426_));
 sky130_fd_sc_hd__and2b_1 _10050_ (.A_N(_04425_),
    .B(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__o21ba_1 _10051_ (.A1(_04395_),
    .A2(_04405_),
    .B1_N(_04393_),
    .X(_04428_));
 sky130_fd_sc_hd__o21ai_1 _10052_ (.A1(_04427_),
    .A2(_04428_),
    .B1(_03867_),
    .Y(_04429_));
 sky130_fd_sc_hd__a21o_1 _10053_ (.A1(_04427_),
    .A2(_04428_),
    .B1(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__o211a_1 _10054_ (.A1(\_185_[21] ),
    .A2(_03870_),
    .B1(_03864_),
    .C1(_04430_),
    .X(_00430_));
 sky130_fd_sc_hd__o221a_1 _10055_ (.A1(\_246_[22] ),
    .A2(_01315_),
    .B1(_04409_),
    .B2(\_243_[22] ),
    .C1(_01497_),
    .X(_04431_));
 sky130_fd_sc_hd__and2_1 _10056_ (.A(\_142_[22] ),
    .B(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__nor2_1 _10057_ (.A(\_142_[22] ),
    .B(_04431_),
    .Y(_04433_));
 sky130_fd_sc_hd__or2_1 _10058_ (.A(_04432_),
    .B(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__a221o_1 _10059_ (.A1(_01244_),
    .A2(_03927_),
    .B1(_03929_),
    .B2(_04156_),
    .C1(_01238_),
    .X(_04435_));
 sky130_fd_sc_hd__nand2_1 _10060_ (.A(_01284_),
    .B(_04005_),
    .Y(_04436_));
 sky130_fd_sc_hd__buf_2 _10061_ (.A(_04078_),
    .X(_04437_));
 sky130_fd_sc_hd__a21oi_1 _10062_ (.A1(_04436_),
    .A2(_04160_),
    .B1(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__nand2_1 _10063_ (.A(_04059_),
    .B(_04438_),
    .Y(_04439_));
 sky130_fd_sc_hd__a32o_1 _10064_ (.A1(_01244_),
    .A2(_04051_),
    .A3(_03903_),
    .B1(_03952_),
    .B2(_03960_),
    .X(_04440_));
 sky130_fd_sc_hd__a2111o_1 _10065_ (.A1(_03873_),
    .A2(_03876_),
    .B1(_04027_),
    .C1(_04303_),
    .D1(_04078_),
    .X(_04441_));
 sky130_fd_sc_hd__o211a_1 _10066_ (.A1(_01238_),
    .A2(_04440_),
    .B1(_04441_),
    .C1(_01232_),
    .X(_04442_));
 sky130_fd_sc_hd__a31o_1 _10067_ (.A1(_04210_),
    .A2(_04435_),
    .A3(_04439_),
    .B1(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__nor2_1 _10068_ (.A(_04434_),
    .B(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__nand2_1 _10069_ (.A(_04434_),
    .B(_04443_),
    .Y(_04445_));
 sky130_fd_sc_hd__and2b_1 _10070_ (.A_N(_04444_),
    .B(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__o21ai_1 _10071_ (.A1(_04411_),
    .A2(_04422_),
    .B1(_04446_),
    .Y(_04447_));
 sky130_fd_sc_hd__or3_1 _10072_ (.A(_04411_),
    .B(_04422_),
    .C(_04446_),
    .X(_04448_));
 sky130_fd_sc_hd__and2_1 _10073_ (.A(_04447_),
    .B(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__or3b_1 _10074_ (.A(_04395_),
    .B(_04425_),
    .C_N(_04426_),
    .X(_04450_));
 sky130_fd_sc_hd__a21oi_2 _10075_ (.A1(_04398_),
    .A2(_04404_),
    .B1(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__o21a_1 _10076_ (.A1(_04393_),
    .A2(_04425_),
    .B1(_04426_),
    .X(_04452_));
 sky130_fd_sc_hd__or2_1 _10077_ (.A(_04451_),
    .B(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__xnor2_1 _10078_ (.A(_04449_),
    .B(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__nand2_1 _10079_ (.A(_03868_),
    .B(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__o211a_1 _10080_ (.A1(\_185_[22] ),
    .A2(_03870_),
    .B1(_03864_),
    .C1(_04455_),
    .X(_00431_));
 sky130_fd_sc_hd__a211o_1 _10081_ (.A1(_03901_),
    .A2(_04160_),
    .B1(_04333_),
    .C1(_03935_),
    .X(_04456_));
 sky130_fd_sc_hd__and4_1 _10082_ (.A(_04060_),
    .B(_03984_),
    .C(_04025_),
    .D(_04418_),
    .X(_04457_));
 sky130_fd_sc_hd__o22a_1 _10083_ (.A1(_01281_),
    .A2(_03934_),
    .B1(_03904_),
    .B2(_03905_),
    .X(_04458_));
 sky130_fd_sc_hd__o21ai_1 _10084_ (.A1(_04075_),
    .A2(_03960_),
    .B1(_04278_),
    .Y(_04459_));
 sky130_fd_sc_hd__o211a_1 _10085_ (.A1(_01238_),
    .A2(_04458_),
    .B1(_04459_),
    .C1(_01232_),
    .X(_04460_));
 sky130_fd_sc_hd__a211o_1 _10086_ (.A1(_04054_),
    .A2(_04456_),
    .B1(_04457_),
    .C1(_04460_),
    .X(_04461_));
 sky130_fd_sc_hd__o221a_1 _10087_ (.A1(\_246_[23] ),
    .A2(_01316_),
    .B1(_04409_),
    .B2(\_243_[23] ),
    .C1(_01499_),
    .X(_04462_));
 sky130_fd_sc_hd__xnor2_1 _10088_ (.A(\_142_[23] ),
    .B(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__xor2_1 _10089_ (.A(_04461_),
    .B(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__nor3_1 _10090_ (.A(_04432_),
    .B(_04444_),
    .C(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__o21a_1 _10091_ (.A1(_04432_),
    .A2(_04444_),
    .B1(_04464_),
    .X(_04466_));
 sky130_fd_sc_hd__nor2_1 _10092_ (.A(_04465_),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__a21boi_1 _10093_ (.A1(_04449_),
    .A2(_04453_),
    .B1_N(_04447_),
    .Y(_04468_));
 sky130_fd_sc_hd__o21ai_1 _10094_ (.A1(_04467_),
    .A2(_04468_),
    .B1(_03867_),
    .Y(_04469_));
 sky130_fd_sc_hd__a21o_1 _10095_ (.A1(_04467_),
    .A2(_04468_),
    .B1(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__o211a_1 _10096_ (.A1(\_185_[23] ),
    .A2(_03870_),
    .B1(_03864_),
    .C1(_04470_),
    .X(_00432_));
 sky130_fd_sc_hd__o221a_1 _10097_ (.A1(\_246_[24] ),
    .A2(_01315_),
    .B1(_04409_),
    .B2(\_243_[24] ),
    .C1(_01501_),
    .X(_04471_));
 sky130_fd_sc_hd__and2_1 _10098_ (.A(\_142_[24] ),
    .B(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__nor2_1 _10099_ (.A(\_142_[24] ),
    .B(_04471_),
    .Y(_04473_));
 sky130_fd_sc_hd__or2_1 _10100_ (.A(_04472_),
    .B(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__nand2_1 _10101_ (.A(_04085_),
    .B(_04177_),
    .Y(_04475_));
 sky130_fd_sc_hd__a2bb2o_1 _10102_ (.A1_N(_01292_),
    .A2_N(_04057_),
    .B1(_04475_),
    .B2(_01238_),
    .X(_04476_));
 sky130_fd_sc_hd__o31a_1 _10103_ (.A1(_03886_),
    .A2(_03976_),
    .A3(_04476_),
    .B1(_01233_),
    .X(_04477_));
 sky130_fd_sc_hd__a311oi_2 _10104_ (.A1(_04436_),
    .A2(_03984_),
    .A3(_04365_),
    .B1(_04318_),
    .C1(_04157_),
    .Y(_04478_));
 sky130_fd_sc_hd__inv_2 _10105_ (.A(_04320_),
    .Y(_04479_));
 sky130_fd_sc_hd__a21oi_1 _10106_ (.A1(_04436_),
    .A2(_04479_),
    .B1(_03906_),
    .Y(_04480_));
 sky130_fd_sc_hd__nor2_1 _10107_ (.A(_04161_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__nor4_1 _10108_ (.A(_04474_),
    .B(_04477_),
    .C(_04478_),
    .D(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__o31a_1 _10109_ (.A1(_04477_),
    .A2(_04478_),
    .A3(_04481_),
    .B1(_04474_),
    .X(_04483_));
 sky130_fd_sc_hd__nor2_1 _10110_ (.A(_04482_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__o2bb2ai_1 _10111_ (.A1_N(\_142_[23] ),
    .A2_N(_04462_),
    .B1(_04463_),
    .B2(_04461_),
    .Y(_04485_));
 sky130_fd_sc_hd__and2_1 _10112_ (.A(_04484_),
    .B(_04485_),
    .X(_04486_));
 sky130_fd_sc_hd__nor2_1 _10113_ (.A(_04484_),
    .B(_04485_),
    .Y(_04487_));
 sky130_fd_sc_hd__nor2_1 _10114_ (.A(_04486_),
    .B(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__o21bai_2 _10115_ (.A1(_04447_),
    .A2(_04465_),
    .B1_N(_04466_),
    .Y(_04489_));
 sky130_fd_sc_hd__a21o_1 _10116_ (.A1(_04449_),
    .A2(_04467_),
    .B1(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__o31a_1 _10117_ (.A1(_04451_),
    .A2(_04452_),
    .A3(_04489_),
    .B1(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__xor2_1 _10118_ (.A(_04488_),
    .B(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__or2_1 _10119_ (.A(\_185_[24] ),
    .B(_03867_),
    .X(_04493_));
 sky130_fd_sc_hd__o211a_1 _10120_ (.A1(_03946_),
    .A2(_04492_),
    .B1(_04493_),
    .C1(_00105_),
    .X(_00433_));
 sky130_fd_sc_hd__o221a_1 _10121_ (.A1(\_246_[25] ),
    .A2(_01316_),
    .B1(_04409_),
    .B2(\_243_[25] ),
    .C1(_01503_),
    .X(_04494_));
 sky130_fd_sc_hd__and2_1 _10122_ (.A(\_142_[25] ),
    .B(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__nor2_1 _10123_ (.A(\_142_[25] ),
    .B(_04494_),
    .Y(_04496_));
 sky130_fd_sc_hd__or2_1 _10124_ (.A(_04495_),
    .B(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__nand2_1 _10125_ (.A(_03887_),
    .B(_03925_),
    .Y(_04498_));
 sky130_fd_sc_hd__o2bb2a_1 _10126_ (.A1_N(_04438_),
    .A2_N(_04498_),
    .B1(_01238_),
    .B2(_04365_),
    .X(_04499_));
 sky130_fd_sc_hd__o21ai_1 _10127_ (.A1(_03979_),
    .A2(_04479_),
    .B1(_01238_),
    .Y(_04500_));
 sky130_fd_sc_hd__o311a_1 _10128_ (.A1(_01238_),
    .A2(_04032_),
    .A3(_04258_),
    .B1(_04500_),
    .C1(_01232_),
    .X(_04501_));
 sky130_fd_sc_hd__inv_2 _10129_ (.A(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__o31a_1 _10130_ (.A1(_01233_),
    .A2(_03978_),
    .A3(_04499_),
    .B1(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__xnor2_1 _10131_ (.A(_04497_),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__o21bai_1 _10132_ (.A1(_04472_),
    .A2(_04482_),
    .B1_N(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__nor3b_1 _10133_ (.A(_04472_),
    .B(_04482_),
    .C_N(_04504_),
    .Y(_04506_));
 sky130_fd_sc_hd__inv_2 _10134_ (.A(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__nand2_1 _10135_ (.A(_04505_),
    .B(_04507_),
    .Y(_04508_));
 sky130_fd_sc_hd__a21o_1 _10136_ (.A1(_04488_),
    .A2(_04491_),
    .B1(_04486_),
    .X(_04509_));
 sky130_fd_sc_hd__xnor2_1 _10137_ (.A(_04508_),
    .B(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__or2_1 _10138_ (.A(\_185_[25] ),
    .B(_03867_),
    .X(_04511_));
 sky130_fd_sc_hd__o211a_1 _10139_ (.A1(_03946_),
    .A2(_04510_),
    .B1(_04511_),
    .C1(_00105_),
    .X(_00434_));
 sky130_fd_sc_hd__nor2_1 _10140_ (.A(_04497_),
    .B(_04503_),
    .Y(_04512_));
 sky130_fd_sc_hd__or2_1 _10141_ (.A(\_243_[26] ),
    .B(_04409_),
    .X(_04513_));
 sky130_fd_sc_hd__o22a_1 _10142_ (.A1(\_246_[26] ),
    .A2(_01316_),
    .B1(_01301_),
    .B2(\_179_[26] ),
    .X(_04514_));
 sky130_fd_sc_hd__and3_1 _10143_ (.A(\_142_[26] ),
    .B(_04513_),
    .C(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__a21oi_1 _10144_ (.A1(_04513_),
    .A2(_04514_),
    .B1(\_142_[26] ),
    .Y(_04516_));
 sky130_fd_sc_hd__or2_1 _10145_ (.A(_04515_),
    .B(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__o21a_1 _10146_ (.A1(_04027_),
    .A2(_03976_),
    .B1(_04103_),
    .X(_04518_));
 sky130_fd_sc_hd__o32a_1 _10147_ (.A1(_01232_),
    .A2(_04333_),
    .A3(_04366_),
    .B1(_04518_),
    .B2(_04362_),
    .X(_04519_));
 sky130_fd_sc_hd__nor2_1 _10148_ (.A(_03935_),
    .B(_04085_),
    .Y(_04520_));
 sky130_fd_sc_hd__a211o_1 _10149_ (.A1(_01281_),
    .A2(_03876_),
    .B1(_04520_),
    .C1(_04210_),
    .X(_04521_));
 sky130_fd_sc_hd__o311a_1 _10150_ (.A1(_01233_),
    .A2(_03903_),
    .A3(_03876_),
    .B1(_04521_),
    .C1(_04437_),
    .X(_04522_));
 sky130_fd_sc_hd__a21o_1 _10151_ (.A1(_01239_),
    .A2(_04519_),
    .B1(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__nor2_1 _10152_ (.A(_04517_),
    .B(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__and2_1 _10153_ (.A(_04517_),
    .B(_04523_),
    .X(_04525_));
 sky130_fd_sc_hd__nor2_1 _10154_ (.A(_04524_),
    .B(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__o21ai_1 _10155_ (.A1(_04495_),
    .A2(_04512_),
    .B1(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__or3_1 _10156_ (.A(_04495_),
    .B(_04512_),
    .C(_04526_),
    .X(_04528_));
 sky130_fd_sc_hd__and2_1 _10157_ (.A(_04527_),
    .B(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__and3_1 _10158_ (.A(_04488_),
    .B(_04505_),
    .C(_04507_),
    .X(_04530_));
 sky130_fd_sc_hd__o311ai_4 _10159_ (.A1(_04451_),
    .A2(_04452_),
    .A3(_04489_),
    .B1(_04490_),
    .C1(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__inv_2 _10160_ (.A(_04486_),
    .Y(_04532_));
 sky130_fd_sc_hd__a21o_1 _10161_ (.A1(_04532_),
    .A2(_04505_),
    .B1(_04506_),
    .X(_04533_));
 sky130_fd_sc_hd__nand2_1 _10162_ (.A(_04531_),
    .B(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__xor2_1 _10163_ (.A(_04529_),
    .B(_04534_),
    .X(_04535_));
 sky130_fd_sc_hd__or2_1 _10164_ (.A(\_185_[26] ),
    .B(_03867_),
    .X(_04536_));
 sky130_fd_sc_hd__o211a_1 _10165_ (.A1(_03946_),
    .A2(_04535_),
    .B1(_04536_),
    .C1(_00105_),
    .X(_00435_));
 sky130_fd_sc_hd__nand2_1 _10166_ (.A(_04529_),
    .B(_04534_),
    .Y(_04537_));
 sky130_fd_sc_hd__o221a_1 _10167_ (.A1(\_246_[27] ),
    .A2(_01316_),
    .B1(_04409_),
    .B2(\_243_[27] ),
    .C1(_01507_),
    .X(_04538_));
 sky130_fd_sc_hd__xnor2_1 _10168_ (.A(\_142_[27] ),
    .B(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__nor2_1 _10169_ (.A(_04103_),
    .B(_03878_),
    .Y(_04540_));
 sky130_fd_sc_hd__or3_1 _10170_ (.A(_04437_),
    .B(_03893_),
    .C(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__nor2_1 _10171_ (.A(_04081_),
    .B(_04010_),
    .Y(_04542_));
 sky130_fd_sc_hd__a211o_1 _10172_ (.A1(_03954_),
    .A2(_04156_),
    .B1(_04542_),
    .C1(_01238_),
    .X(_04543_));
 sky130_fd_sc_hd__nand2_1 _10173_ (.A(_04437_),
    .B(_04108_),
    .Y(_04544_));
 sky130_fd_sc_hd__o221a_1 _10174_ (.A1(_03899_),
    .A2(_04215_),
    .B1(_04544_),
    .B2(_03925_),
    .C1(_01233_),
    .X(_04545_));
 sky130_fd_sc_hd__a31o_1 _10175_ (.A1(_04210_),
    .A2(_04541_),
    .A3(_04543_),
    .B1(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__xnor2_1 _10176_ (.A(_04539_),
    .B(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__nor3b_1 _10177_ (.A(_04515_),
    .B(_04524_),
    .C_N(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__o21ba_1 _10178_ (.A1(_04515_),
    .A2(_04524_),
    .B1_N(_04547_),
    .X(_04549_));
 sky130_fd_sc_hd__nor2_1 _10179_ (.A(_04548_),
    .B(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__and3_1 _10180_ (.A(_04527_),
    .B(_04537_),
    .C(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__a21oi_1 _10181_ (.A1(_04527_),
    .A2(_04537_),
    .B1(_04550_),
    .Y(_04552_));
 sky130_fd_sc_hd__or3_1 _10182_ (.A(_03945_),
    .B(_04551_),
    .C(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__o211a_1 _10183_ (.A1(\_185_[27] ),
    .A2(_03870_),
    .B1(_03864_),
    .C1(_04553_),
    .X(_00436_));
 sky130_fd_sc_hd__nand2_1 _10184_ (.A(_04529_),
    .B(_04550_),
    .Y(_04554_));
 sky130_fd_sc_hd__o21ba_1 _10185_ (.A1(_04527_),
    .A2(_04548_),
    .B1_N(_04549_),
    .X(_04555_));
 sky130_fd_sc_hd__and2_1 _10186_ (.A(_04533_),
    .B(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__o221a_1 _10187_ (.A1(\_246_[28] ),
    .A2(_01316_),
    .B1(_04409_),
    .B2(\_243_[28] ),
    .C1(_01511_),
    .X(_04557_));
 sky130_fd_sc_hd__and2_1 _10188_ (.A(\_142_[28] ),
    .B(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__nor2_1 _10189_ (.A(\_142_[28] ),
    .B(_04557_),
    .Y(_04559_));
 sky130_fd_sc_hd__or2_1 _10190_ (.A(_04558_),
    .B(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__o32a_1 _10191_ (.A1(_04437_),
    .A2(_03952_),
    .A3(_04026_),
    .B1(_04540_),
    .B2(_03894_),
    .X(_04561_));
 sky130_fd_sc_hd__o21a_1 _10192_ (.A1(_04303_),
    .A2(_04233_),
    .B1(_04437_),
    .X(_04562_));
 sky130_fd_sc_hd__a41o_1 _10193_ (.A1(_01239_),
    .A2(_03890_),
    .A3(_03888_),
    .A4(_03938_),
    .B1(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__mux2_1 _10194_ (.A0(_04561_),
    .A1(_04563_),
    .S(_01233_),
    .X(_04564_));
 sky130_fd_sc_hd__xnor2_1 _10195_ (.A(_04560_),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__o2bb2a_1 _10196_ (.A1_N(\_142_[27] ),
    .A2_N(_04538_),
    .B1(_04539_),
    .B2(_04546_),
    .X(_04566_));
 sky130_fd_sc_hd__xnor2_1 _10197_ (.A(_04565_),
    .B(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__a221oi_4 _10198_ (.A1(_04554_),
    .A2(_04555_),
    .B1(_04556_),
    .B2(_04531_),
    .C1(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__a22o_1 _10199_ (.A1(_04554_),
    .A2(_04555_),
    .B1(_04556_),
    .B2(_04531_),
    .X(_04569_));
 sky130_fd_sc_hd__and2_1 _10200_ (.A(_04567_),
    .B(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__o21ai_1 _10201_ (.A1(_04568_),
    .A2(_04570_),
    .B1(_03868_),
    .Y(_04571_));
 sky130_fd_sc_hd__o211a_1 _10202_ (.A1(\_185_[28] ),
    .A2(_03870_),
    .B1(_03864_),
    .C1(_04571_),
    .X(_00437_));
 sky130_fd_sc_hd__nor2_1 _10203_ (.A(_04565_),
    .B(_04566_),
    .Y(_04572_));
 sky130_fd_sc_hd__nor2_1 _10204_ (.A(_04560_),
    .B(_04564_),
    .Y(_04573_));
 sky130_fd_sc_hd__or3_1 _10205_ (.A(_04437_),
    .B(_04158_),
    .C(_04360_),
    .X(_04574_));
 sky130_fd_sc_hd__o31a_1 _10206_ (.A1(_01239_),
    .A2(_04163_),
    .A3(_04416_),
    .B1(_04210_),
    .X(_04575_));
 sky130_fd_sc_hd__a21o_1 _10207_ (.A1(_03890_),
    .A2(_03927_),
    .B1(_01244_),
    .X(_04576_));
 sky130_fd_sc_hd__o211a_1 _10208_ (.A1(_04303_),
    .A2(_04085_),
    .B1(_04576_),
    .C1(_01239_),
    .X(_04577_));
 sky130_fd_sc_hd__o21ai_1 _10209_ (.A1(_04303_),
    .A2(_04103_),
    .B1(_04135_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand2_1 _10210_ (.A(_01233_),
    .B(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__o2bb2a_1 _10211_ (.A1_N(_04574_),
    .A2_N(_04575_),
    .B1(_04577_),
    .B2(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__o221a_1 _10212_ (.A1(\_246_[29] ),
    .A2(_01316_),
    .B1(_04409_),
    .B2(\_243_[29] ),
    .C1(_01513_),
    .X(_04581_));
 sky130_fd_sc_hd__and2_1 _10213_ (.A(\_142_[29] ),
    .B(_04581_),
    .X(_04582_));
 sky130_fd_sc_hd__nor2_1 _10214_ (.A(\_142_[29] ),
    .B(_04581_),
    .Y(_04583_));
 sky130_fd_sc_hd__nor2_1 _10215_ (.A(_04582_),
    .B(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__and2_1 _10216_ (.A(_04580_),
    .B(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__nor2_1 _10217_ (.A(_04580_),
    .B(_04584_),
    .Y(_04586_));
 sky130_fd_sc_hd__or2_1 _10218_ (.A(_04585_),
    .B(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__o21ba_1 _10219_ (.A1(_04558_),
    .A2(_04573_),
    .B1_N(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__or3b_1 _10220_ (.A(_04558_),
    .B(_04573_),
    .C_N(_04587_),
    .X(_04589_));
 sky130_fd_sc_hd__or2b_1 _10221_ (.A(_04588_),
    .B_N(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__nor3_1 _10222_ (.A(_04572_),
    .B(_04568_),
    .C(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__o21a_1 _10223_ (.A1(_04572_),
    .A2(_04568_),
    .B1(_04590_),
    .X(_04592_));
 sky130_fd_sc_hd__or3_1 _10224_ (.A(_03945_),
    .B(_04591_),
    .C(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__o211a_1 _10225_ (.A1(\_185_[29] ),
    .A2(_03870_),
    .B1(_03864_),
    .C1(_04593_),
    .X(_00438_));
 sky130_fd_sc_hd__a32o_1 _10226_ (.A1(_03896_),
    .A2(_04132_),
    .A3(_03984_),
    .B1(_03878_),
    .B2(_01244_),
    .X(_04594_));
 sky130_fd_sc_hd__nor2_1 _10227_ (.A(_01239_),
    .B(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__nor2_1 _10228_ (.A(_04164_),
    .B(_04386_),
    .Y(_04596_));
 sky130_fd_sc_hd__o211a_1 _10229_ (.A1(_03950_),
    .A2(_04363_),
    .B1(_03890_),
    .C1(_04437_),
    .X(_04597_));
 sky130_fd_sc_hd__o211a_1 _10230_ (.A1(_01285_),
    .A2(_04107_),
    .B1(_04385_),
    .C1(_01239_),
    .X(_04598_));
 sky130_fd_sc_hd__or3_1 _10231_ (.A(_04210_),
    .B(_04597_),
    .C(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__o31a_1 _10232_ (.A1(_01233_),
    .A2(_04595_),
    .A3(_04596_),
    .B1(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__o221a_2 _10233_ (.A1(\_246_[30] ),
    .A2(_01316_),
    .B1(_04409_),
    .B2(\_243_[30] ),
    .C1(_01516_),
    .X(_04601_));
 sky130_fd_sc_hd__xor2_1 _10234_ (.A(\_142_[30] ),
    .B(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__xnor2_1 _10235_ (.A(_04600_),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__o21ba_1 _10236_ (.A1(_04582_),
    .A2(_04585_),
    .B1_N(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__or3b_1 _10237_ (.A(_04582_),
    .B(_04585_),
    .C_N(_04603_),
    .X(_04605_));
 sky130_fd_sc_hd__and2b_1 _10238_ (.A_N(_04604_),
    .B(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__o31a_1 _10239_ (.A1(_04572_),
    .A2(_04568_),
    .A3(_04588_),
    .B1(_04589_),
    .X(_04607_));
 sky130_fd_sc_hd__xor2_1 _10240_ (.A(_04606_),
    .B(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__or2_1 _10241_ (.A(\_185_[30] ),
    .B(_03867_),
    .X(_04609_));
 sky130_fd_sc_hd__o211a_1 _10242_ (.A1(_03946_),
    .A2(_04608_),
    .B1(_04609_),
    .C1(_00105_),
    .X(_00439_));
 sky130_fd_sc_hd__a21oi_1 _10243_ (.A1(_04605_),
    .A2(_04607_),
    .B1(_04604_),
    .Y(_04610_));
 sky130_fd_sc_hd__mux2_1 _10244_ (.A0(\_246_[31] ),
    .A1(\_243_[31] ),
    .S(_01316_),
    .X(_04611_));
 sky130_fd_sc_hd__a21oi_2 _10245_ (.A1(_01353_),
    .A2(_04611_),
    .B1(_01521_),
    .Y(_04612_));
 sky130_fd_sc_hd__a22o_1 _10246_ (.A1(\_142_[30] ),
    .A2(_04601_),
    .B1(_04602_),
    .B2(_04600_),
    .X(_04613_));
 sky130_fd_sc_hd__or3_1 _10247_ (.A(_04055_),
    .B(_04077_),
    .C(_04361_),
    .X(_04614_));
 sky130_fd_sc_hd__or3b_1 _10248_ (.A(_04132_),
    .B(_04437_),
    .C_N(_03950_),
    .X(_04615_));
 sky130_fd_sc_hd__a211o_1 _10249_ (.A1(_01244_),
    .A2(_01285_),
    .B1(_03952_),
    .C1(_01239_),
    .X(_04616_));
 sky130_fd_sc_hd__o211a_1 _10250_ (.A1(_04437_),
    .A2(_04107_),
    .B1(_04616_),
    .C1(_01233_),
    .X(_04617_));
 sky130_fd_sc_hd__a31o_1 _10251_ (.A1(_04210_),
    .A2(_04614_),
    .A3(_04615_),
    .B1(_04617_),
    .X(_04618_));
 sky130_fd_sc_hd__xnor2_1 _10252_ (.A(\_142_[31] ),
    .B(_04618_),
    .Y(_04619_));
 sky130_fd_sc_hd__xnor2_1 _10253_ (.A(_04613_),
    .B(_04619_),
    .Y(_04620_));
 sky130_fd_sc_hd__xnor2_1 _10254_ (.A(_04612_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__xnor2_1 _10255_ (.A(_04610_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__o21ai_1 _10256_ (.A1(\_185_[31] ),
    .A2(_03868_),
    .B1(_03864_),
    .Y(_04623_));
 sky130_fd_sc_hd__a21oi_1 _10257_ (.A1(_03870_),
    .A2(_04622_),
    .B1(_04623_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand2_1 _10258_ (.A(_01272_),
    .B(_01349_),
    .Y(_04624_));
 sky130_fd_sc_hd__nor3_4 _10259_ (.A(_01305_),
    .B(_01338_),
    .C(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__nand2_1 _10260_ (.A(_01212_),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__buf_4 _10261_ (.A(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__clkbuf_4 _10262_ (.A(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__buf_4 _10263_ (.A(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__buf_4 _10264_ (.A(_04625_),
    .X(_04630_));
 sky130_fd_sc_hd__buf_4 _10265_ (.A(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__a31o_1 _10266_ (.A1(\_182_[0] ),
    .A2(_01218_),
    .A3(_04631_),
    .B1(_03309_),
    .X(_04632_));
 sky130_fd_sc_hd__a21o_1 _10267_ (.A1(\_179_[0] ),
    .A2(_04629_),
    .B1(_04632_),
    .X(_00441_));
 sky130_fd_sc_hd__buf_4 _10268_ (.A(_04626_),
    .X(_04633_));
 sky130_fd_sc_hd__clkbuf_4 _10269_ (.A(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__or3_2 _10270_ (.A(_01305_),
    .B(_01338_),
    .C(_04624_),
    .X(_04635_));
 sky130_fd_sc_hd__buf_4 _10271_ (.A(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__nor2_4 _10272_ (.A(_01214_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__buf_4 _10273_ (.A(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__or2_1 _10274_ (.A(\_179_[1] ),
    .B(_04638_),
    .X(_04639_));
 sky130_fd_sc_hd__o211a_1 _10275_ (.A1(\_182_[1] ),
    .A2(_04634_),
    .B1(_04639_),
    .C1(_00105_),
    .X(_00442_));
 sky130_fd_sc_hd__or2_1 _10276_ (.A(\_179_[2] ),
    .B(_04638_),
    .X(_04640_));
 sky130_fd_sc_hd__o211a_1 _10277_ (.A1(\_182_[2] ),
    .A2(_04634_),
    .B1(_04640_),
    .C1(_00105_),
    .X(_00443_));
 sky130_fd_sc_hd__a31o_1 _10278_ (.A1(\_182_[3] ),
    .A2(_01218_),
    .A3(_04631_),
    .B1(_03309_),
    .X(_04641_));
 sky130_fd_sc_hd__a21o_1 _10279_ (.A1(\_179_[3] ),
    .A2(_04629_),
    .B1(_04641_),
    .X(_00444_));
 sky130_fd_sc_hd__clkbuf_4 _10280_ (.A(_04630_),
    .X(_04642_));
 sky130_fd_sc_hd__a31o_1 _10281_ (.A1(\_182_[4] ),
    .A2(_01218_),
    .A3(_04642_),
    .B1(_03309_),
    .X(_04643_));
 sky130_fd_sc_hd__a21o_1 _10282_ (.A1(\_179_[4] ),
    .A2(_04629_),
    .B1(_04643_),
    .X(_00445_));
 sky130_fd_sc_hd__or2_1 _10283_ (.A(\_179_[5] ),
    .B(_04638_),
    .X(_04644_));
 sky130_fd_sc_hd__o211a_1 _10284_ (.A1(\_182_[5] ),
    .A2(_04634_),
    .B1(_04644_),
    .C1(_00105_),
    .X(_00446_));
 sky130_fd_sc_hd__or2_1 _10285_ (.A(\_179_[6] ),
    .B(_04638_),
    .X(_04645_));
 sky130_fd_sc_hd__o211a_1 _10286_ (.A1(\_182_[6] ),
    .A2(_04634_),
    .B1(_04645_),
    .C1(_00105_),
    .X(_00447_));
 sky130_fd_sc_hd__clkbuf_4 _10287_ (.A(_04637_),
    .X(_04646_));
 sky130_fd_sc_hd__or2_1 _10288_ (.A(\_179_[7] ),
    .B(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__clkbuf_8 _10289_ (.A(_01423_),
    .X(_04648_));
 sky130_fd_sc_hd__clkbuf_4 _10290_ (.A(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__o211a_1 _10291_ (.A1(\_182_[7] ),
    .A2(_04634_),
    .B1(_04647_),
    .C1(_04649_),
    .X(_00448_));
 sky130_fd_sc_hd__clkbuf_4 _10292_ (.A(_01417_),
    .X(_04650_));
 sky130_fd_sc_hd__a31o_1 _10293_ (.A1(\_182_[8] ),
    .A2(_01218_),
    .A3(_04642_),
    .B1(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__a21o_1 _10294_ (.A1(\_179_[8] ),
    .A2(_04629_),
    .B1(_04651_),
    .X(_00449_));
 sky130_fd_sc_hd__or2_1 _10295_ (.A(\_179_[9] ),
    .B(_04646_),
    .X(_04652_));
 sky130_fd_sc_hd__o211a_1 _10296_ (.A1(\_182_[9] ),
    .A2(_04634_),
    .B1(_04652_),
    .C1(_04649_),
    .X(_00450_));
 sky130_fd_sc_hd__a31o_1 _10297_ (.A1(\_182_[10] ),
    .A2(_01218_),
    .A3(_04642_),
    .B1(_04650_),
    .X(_04653_));
 sky130_fd_sc_hd__a21o_1 _10298_ (.A1(\_179_[10] ),
    .A2(_04629_),
    .B1(_04653_),
    .X(_00451_));
 sky130_fd_sc_hd__clkbuf_4 _10299_ (.A(_01217_),
    .X(_04654_));
 sky130_fd_sc_hd__a31o_1 _10300_ (.A1(\_182_[11] ),
    .A2(_04654_),
    .A3(_04642_),
    .B1(_04650_),
    .X(_04655_));
 sky130_fd_sc_hd__a21o_1 _10301_ (.A1(\_179_[11] ),
    .A2(_04629_),
    .B1(_04655_),
    .X(_00452_));
 sky130_fd_sc_hd__or2_1 _10302_ (.A(\_179_[12] ),
    .B(_04646_),
    .X(_04656_));
 sky130_fd_sc_hd__o211a_1 _10303_ (.A1(\_182_[12] ),
    .A2(_04634_),
    .B1(_04656_),
    .C1(_04649_),
    .X(_00453_));
 sky130_fd_sc_hd__or2_1 _10304_ (.A(\_179_[13] ),
    .B(_04646_),
    .X(_04657_));
 sky130_fd_sc_hd__o211a_1 _10305_ (.A1(\_182_[13] ),
    .A2(_04634_),
    .B1(_04657_),
    .C1(_04649_),
    .X(_00454_));
 sky130_fd_sc_hd__clkbuf_4 _10306_ (.A(_04633_),
    .X(_04658_));
 sky130_fd_sc_hd__a31o_1 _10307_ (.A1(\_182_[14] ),
    .A2(_04654_),
    .A3(_04642_),
    .B1(_04650_),
    .X(_04659_));
 sky130_fd_sc_hd__a21o_1 _10308_ (.A1(\_179_[14] ),
    .A2(_04658_),
    .B1(_04659_),
    .X(_00455_));
 sky130_fd_sc_hd__a31o_1 _10309_ (.A1(\_182_[15] ),
    .A2(_04654_),
    .A3(_04642_),
    .B1(_04650_),
    .X(_04660_));
 sky130_fd_sc_hd__a21o_1 _10310_ (.A1(\_179_[15] ),
    .A2(_04658_),
    .B1(_04660_),
    .X(_00456_));
 sky130_fd_sc_hd__or2_1 _10311_ (.A(\_179_[16] ),
    .B(_04646_),
    .X(_04661_));
 sky130_fd_sc_hd__o211a_1 _10312_ (.A1(\_182_[16] ),
    .A2(_04634_),
    .B1(_04661_),
    .C1(_04649_),
    .X(_00457_));
 sky130_fd_sc_hd__or2_1 _10313_ (.A(\_179_[17] ),
    .B(_04646_),
    .X(_04662_));
 sky130_fd_sc_hd__o211a_1 _10314_ (.A1(\_182_[17] ),
    .A2(_04634_),
    .B1(_04662_),
    .C1(_04649_),
    .X(_00458_));
 sky130_fd_sc_hd__clkbuf_4 _10315_ (.A(_04633_),
    .X(_04663_));
 sky130_fd_sc_hd__or2_1 _10316_ (.A(\_179_[18] ),
    .B(_04646_),
    .X(_04664_));
 sky130_fd_sc_hd__o211a_1 _10317_ (.A1(\_182_[18] ),
    .A2(_04663_),
    .B1(_04664_),
    .C1(_04649_),
    .X(_00459_));
 sky130_fd_sc_hd__or2_1 _10318_ (.A(\_179_[19] ),
    .B(_04646_),
    .X(_04665_));
 sky130_fd_sc_hd__o211a_1 _10319_ (.A1(\_182_[19] ),
    .A2(_04663_),
    .B1(_04665_),
    .C1(_04649_),
    .X(_00460_));
 sky130_fd_sc_hd__or2_1 _10320_ (.A(\_179_[20] ),
    .B(_04646_),
    .X(_04666_));
 sky130_fd_sc_hd__o211a_1 _10321_ (.A1(\_182_[20] ),
    .A2(_04663_),
    .B1(_04666_),
    .C1(_04649_),
    .X(_00461_));
 sky130_fd_sc_hd__a31o_1 _10322_ (.A1(\_182_[21] ),
    .A2(_04654_),
    .A3(_04642_),
    .B1(_04650_),
    .X(_04667_));
 sky130_fd_sc_hd__a21o_1 _10323_ (.A1(\_179_[21] ),
    .A2(_04658_),
    .B1(_04667_),
    .X(_00462_));
 sky130_fd_sc_hd__a31o_1 _10324_ (.A1(\_182_[22] ),
    .A2(_04654_),
    .A3(_04642_),
    .B1(_04650_),
    .X(_04668_));
 sky130_fd_sc_hd__a21o_1 _10325_ (.A1(\_179_[22] ),
    .A2(_04658_),
    .B1(_04668_),
    .X(_00463_));
 sky130_fd_sc_hd__a31o_1 _10326_ (.A1(\_182_[23] ),
    .A2(_04654_),
    .A3(_04642_),
    .B1(_04650_),
    .X(_04669_));
 sky130_fd_sc_hd__a21o_1 _10327_ (.A1(\_179_[23] ),
    .A2(_04658_),
    .B1(_04669_),
    .X(_00464_));
 sky130_fd_sc_hd__a31o_1 _10328_ (.A1(\_182_[24] ),
    .A2(_04654_),
    .A3(_04642_),
    .B1(_04650_),
    .X(_04670_));
 sky130_fd_sc_hd__a21o_1 _10329_ (.A1(\_179_[24] ),
    .A2(_04658_),
    .B1(_04670_),
    .X(_00465_));
 sky130_fd_sc_hd__clkbuf_4 _10330_ (.A(_04630_),
    .X(_04671_));
 sky130_fd_sc_hd__a31o_1 _10331_ (.A1(\_182_[25] ),
    .A2(_04654_),
    .A3(_04671_),
    .B1(_04650_),
    .X(_04672_));
 sky130_fd_sc_hd__a21o_1 _10332_ (.A1(\_179_[25] ),
    .A2(_04658_),
    .B1(_04672_),
    .X(_00466_));
 sky130_fd_sc_hd__or2_1 _10333_ (.A(\_179_[26] ),
    .B(_04646_),
    .X(_04673_));
 sky130_fd_sc_hd__o211a_1 _10334_ (.A1(\_182_[26] ),
    .A2(_04663_),
    .B1(_04673_),
    .C1(_04649_),
    .X(_00467_));
 sky130_fd_sc_hd__a31o_1 _10335_ (.A1(\_182_[27] ),
    .A2(_04654_),
    .A3(_04671_),
    .B1(_01710_),
    .X(_04674_));
 sky130_fd_sc_hd__a21o_1 _10336_ (.A1(\_179_[27] ),
    .A2(_04658_),
    .B1(_04674_),
    .X(_00468_));
 sky130_fd_sc_hd__a31o_1 _10337_ (.A1(\_182_[28] ),
    .A2(_04654_),
    .A3(_04671_),
    .B1(_01710_),
    .X(_04675_));
 sky130_fd_sc_hd__a21o_1 _10338_ (.A1(\_179_[28] ),
    .A2(_04658_),
    .B1(_04675_),
    .X(_00469_));
 sky130_fd_sc_hd__or2_1 _10339_ (.A(\_179_[29] ),
    .B(_04637_),
    .X(_04676_));
 sky130_fd_sc_hd__clkbuf_4 _10340_ (.A(_01424_),
    .X(_04677_));
 sky130_fd_sc_hd__o211a_1 _10341_ (.A1(\_182_[29] ),
    .A2(_04663_),
    .B1(_04676_),
    .C1(_04677_),
    .X(_00470_));
 sky130_fd_sc_hd__buf_4 _10342_ (.A(_01217_),
    .X(_04678_));
 sky130_fd_sc_hd__a31o_1 _10343_ (.A1(\_182_[30] ),
    .A2(_04678_),
    .A3(_04671_),
    .B1(_01710_),
    .X(_04679_));
 sky130_fd_sc_hd__a21o_1 _10344_ (.A1(\_179_[30] ),
    .A2(_04658_),
    .B1(_04679_),
    .X(_00471_));
 sky130_fd_sc_hd__or2_1 _10345_ (.A(\_179_[31] ),
    .B(_04637_),
    .X(_04680_));
 sky130_fd_sc_hd__o211a_1 _10346_ (.A1(\_182_[31] ),
    .A2(_04663_),
    .B1(_04680_),
    .C1(_04677_),
    .X(_00472_));
 sky130_fd_sc_hd__buf_4 _10347_ (.A(_04635_),
    .X(_04681_));
 sky130_fd_sc_hd__clkbuf_4 _10348_ (.A(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__buf_4 _10349_ (.A(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__clkbuf_4 _10350_ (.A(_01225_),
    .X(_04684_));
 sky130_fd_sc_hd__buf_2 _10351_ (.A(_04625_),
    .X(_04685_));
 sky130_fd_sc_hd__clkbuf_4 _10352_ (.A(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__or2_1 _10353_ (.A(\_182_[0] ),
    .B(_01217_),
    .X(_04687_));
 sky130_fd_sc_hd__o211a_1 _10354_ (.A1(\_179_[0] ),
    .A2(_04684_),
    .B1(_04686_),
    .C1(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__a211o_1 _10355_ (.A1(\_176_[0] ),
    .A2(_04683_),
    .B1(_04688_),
    .C1(_01419_),
    .X(_00473_));
 sky130_fd_sc_hd__or2_1 _10356_ (.A(\_182_[1] ),
    .B(_01217_),
    .X(_04689_));
 sky130_fd_sc_hd__o211a_1 _10357_ (.A1(\_179_[1] ),
    .A2(_04684_),
    .B1(_04686_),
    .C1(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__a211o_1 _10358_ (.A1(\_176_[1] ),
    .A2(_04683_),
    .B1(_04690_),
    .C1(_01419_),
    .X(_00474_));
 sky130_fd_sc_hd__clkbuf_8 _10359_ (.A(_04686_),
    .X(_04691_));
 sky130_fd_sc_hd__buf_4 _10360_ (.A(_04636_),
    .X(_04692_));
 sky130_fd_sc_hd__buf_4 _10361_ (.A(_01214_),
    .X(_04693_));
 sky130_fd_sc_hd__mux2_1 _10362_ (.A0(\_179_[2] ),
    .A1(\_182_[2] ),
    .S(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__or2_1 _10363_ (.A(_04692_),
    .B(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__o211a_1 _10364_ (.A1(\_176_[2] ),
    .A2(_04691_),
    .B1(_04695_),
    .C1(_04677_),
    .X(_00475_));
 sky130_fd_sc_hd__buf_2 _10365_ (.A(_01216_),
    .X(_04696_));
 sky130_fd_sc_hd__or2_1 _10366_ (.A(\_182_[3] ),
    .B(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__o211a_1 _10367_ (.A1(\_179_[3] ),
    .A2(_04684_),
    .B1(_04686_),
    .C1(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__a211o_1 _10368_ (.A1(\_176_[3] ),
    .A2(_04683_),
    .B1(_04698_),
    .C1(_01419_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _10369_ (.A0(\_179_[4] ),
    .A1(\_182_[4] ),
    .S(_04693_),
    .X(_04699_));
 sky130_fd_sc_hd__or2_1 _10370_ (.A(_04692_),
    .B(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__o211a_1 _10371_ (.A1(\_176_[4] ),
    .A2(_04691_),
    .B1(_04700_),
    .C1(_04677_),
    .X(_00477_));
 sky130_fd_sc_hd__or2_1 _10372_ (.A(\_182_[5] ),
    .B(_04696_),
    .X(_04701_));
 sky130_fd_sc_hd__o211a_1 _10373_ (.A1(\_179_[5] ),
    .A2(_04684_),
    .B1(_04686_),
    .C1(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__a211o_1 _10374_ (.A1(\_176_[5] ),
    .A2(_04683_),
    .B1(_04702_),
    .C1(_01419_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _10375_ (.A0(\_179_[6] ),
    .A1(\_182_[6] ),
    .S(_04693_),
    .X(_04703_));
 sky130_fd_sc_hd__or2_1 _10376_ (.A(_04692_),
    .B(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__o211a_1 _10377_ (.A1(\_176_[6] ),
    .A2(_04691_),
    .B1(_04704_),
    .C1(_04677_),
    .X(_00479_));
 sky130_fd_sc_hd__clkbuf_4 _10378_ (.A(_04685_),
    .X(_04705_));
 sky130_fd_sc_hd__or2_1 _10379_ (.A(\_182_[7] ),
    .B(_04696_),
    .X(_04706_));
 sky130_fd_sc_hd__o211a_1 _10380_ (.A1(\_179_[7] ),
    .A2(_04684_),
    .B1(_04705_),
    .C1(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__a211o_1 _10381_ (.A1(\_176_[7] ),
    .A2(_04683_),
    .B1(_04707_),
    .C1(_01419_),
    .X(_00480_));
 sky130_fd_sc_hd__or2_1 _10382_ (.A(\_182_[8] ),
    .B(_04696_),
    .X(_04708_));
 sky130_fd_sc_hd__o211a_1 _10383_ (.A1(\_179_[8] ),
    .A2(_04684_),
    .B1(_04705_),
    .C1(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__a211o_1 _10384_ (.A1(\_176_[8] ),
    .A2(_04683_),
    .B1(_04709_),
    .C1(_01419_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _10385_ (.A0(\_179_[9] ),
    .A1(\_182_[9] ),
    .S(_04693_),
    .X(_04710_));
 sky130_fd_sc_hd__or2_1 _10386_ (.A(_04692_),
    .B(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__o211a_1 _10387_ (.A1(\_176_[9] ),
    .A2(_04691_),
    .B1(_04711_),
    .C1(_04677_),
    .X(_00482_));
 sky130_fd_sc_hd__buf_2 _10388_ (.A(_04681_),
    .X(_04712_));
 sky130_fd_sc_hd__mux2_1 _10389_ (.A0(\_179_[10] ),
    .A1(\_182_[10] ),
    .S(_04693_),
    .X(_04713_));
 sky130_fd_sc_hd__or2_1 _10390_ (.A(_04712_),
    .B(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__o211a_1 _10391_ (.A1(\_176_[10] ),
    .A2(_04691_),
    .B1(_04714_),
    .C1(_04677_),
    .X(_00483_));
 sky130_fd_sc_hd__or2_1 _10392_ (.A(\_182_[11] ),
    .B(_04696_),
    .X(_04715_));
 sky130_fd_sc_hd__o211a_1 _10393_ (.A1(\_179_[11] ),
    .A2(_04684_),
    .B1(_04705_),
    .C1(_04715_),
    .X(_04716_));
 sky130_fd_sc_hd__a211o_1 _10394_ (.A1(\_176_[11] ),
    .A2(_04683_),
    .B1(_04716_),
    .C1(_01419_),
    .X(_00484_));
 sky130_fd_sc_hd__or2_1 _10395_ (.A(\_182_[12] ),
    .B(_04696_),
    .X(_04717_));
 sky130_fd_sc_hd__o211a_1 _10396_ (.A1(\_179_[12] ),
    .A2(_04684_),
    .B1(_04705_),
    .C1(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__a211o_1 _10397_ (.A1(\_176_[12] ),
    .A2(_04683_),
    .B1(_04718_),
    .C1(_01419_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _10398_ (.A0(\_179_[13] ),
    .A1(\_182_[13] ),
    .S(_04693_),
    .X(_04719_));
 sky130_fd_sc_hd__or2_1 _10399_ (.A(_04712_),
    .B(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__o211a_1 _10400_ (.A1(\_176_[13] ),
    .A2(_04691_),
    .B1(_04720_),
    .C1(_04677_),
    .X(_00486_));
 sky130_fd_sc_hd__buf_2 _10401_ (.A(_01225_),
    .X(_04721_));
 sky130_fd_sc_hd__or2_1 _10402_ (.A(\_182_[14] ),
    .B(_04696_),
    .X(_04722_));
 sky130_fd_sc_hd__o211a_1 _10403_ (.A1(\_179_[14] ),
    .A2(_04721_),
    .B1(_04705_),
    .C1(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__a211o_1 _10404_ (.A1(\_176_[14] ),
    .A2(_04683_),
    .B1(_04723_),
    .C1(_01419_),
    .X(_00487_));
 sky130_fd_sc_hd__buf_4 _10405_ (.A(_04681_),
    .X(_04724_));
 sky130_fd_sc_hd__buf_2 _10406_ (.A(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__or2_1 _10407_ (.A(\_182_[15] ),
    .B(_04696_),
    .X(_04726_));
 sky130_fd_sc_hd__o211a_1 _10408_ (.A1(\_179_[15] ),
    .A2(_04721_),
    .B1(_04705_),
    .C1(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__clkbuf_4 _10409_ (.A(_01418_),
    .X(_04728_));
 sky130_fd_sc_hd__a211o_1 _10410_ (.A1(\_176_[15] ),
    .A2(_04725_),
    .B1(_04727_),
    .C1(_04728_),
    .X(_00488_));
 sky130_fd_sc_hd__or2_1 _10411_ (.A(\_182_[16] ),
    .B(_04696_),
    .X(_04729_));
 sky130_fd_sc_hd__o211a_1 _10412_ (.A1(\_179_[16] ),
    .A2(_04721_),
    .B1(_04705_),
    .C1(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__a211o_1 _10413_ (.A1(\_176_[16] ),
    .A2(_04725_),
    .B1(_04730_),
    .C1(_04728_),
    .X(_00489_));
 sky130_fd_sc_hd__or2_1 _10414_ (.A(\_182_[17] ),
    .B(_04696_),
    .X(_04731_));
 sky130_fd_sc_hd__o211a_1 _10415_ (.A1(\_179_[17] ),
    .A2(_04721_),
    .B1(_04705_),
    .C1(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__a211o_1 _10416_ (.A1(\_176_[17] ),
    .A2(_04725_),
    .B1(_04732_),
    .C1(_04728_),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _10417_ (.A0(\_179_[18] ),
    .A1(\_182_[18] ),
    .S(_04693_),
    .X(_04733_));
 sky130_fd_sc_hd__or2_1 _10418_ (.A(_04712_),
    .B(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__o211a_1 _10419_ (.A1(\_176_[18] ),
    .A2(_04691_),
    .B1(_04734_),
    .C1(_04677_),
    .X(_00491_));
 sky130_fd_sc_hd__clkbuf_4 _10420_ (.A(_04671_),
    .X(_04735_));
 sky130_fd_sc_hd__mux2_1 _10421_ (.A0(\_179_[19] ),
    .A1(\_182_[19] ),
    .S(_04693_),
    .X(_04736_));
 sky130_fd_sc_hd__or2_1 _10422_ (.A(_04712_),
    .B(_04736_),
    .X(_04737_));
 sky130_fd_sc_hd__o211a_1 _10423_ (.A1(\_176_[19] ),
    .A2(_04735_),
    .B1(_04737_),
    .C1(_04677_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _10424_ (.A0(\_179_[20] ),
    .A1(\_182_[20] ),
    .S(_04693_),
    .X(_04738_));
 sky130_fd_sc_hd__or2_1 _10425_ (.A(_04712_),
    .B(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__clkbuf_4 _10426_ (.A(_01424_),
    .X(_04740_));
 sky130_fd_sc_hd__o211a_1 _10427_ (.A1(\_176_[20] ),
    .A2(_04735_),
    .B1(_04739_),
    .C1(_04740_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _10428_ (.A0(\_179_[21] ),
    .A1(\_182_[21] ),
    .S(_04693_),
    .X(_04741_));
 sky130_fd_sc_hd__or2_1 _10429_ (.A(_04712_),
    .B(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__o211a_1 _10430_ (.A1(\_176_[21] ),
    .A2(_04735_),
    .B1(_04742_),
    .C1(_04740_),
    .X(_00494_));
 sky130_fd_sc_hd__buf_4 _10431_ (.A(_01214_),
    .X(_04743_));
 sky130_fd_sc_hd__mux2_1 _10432_ (.A0(\_179_[22] ),
    .A1(\_182_[22] ),
    .S(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__or2_1 _10433_ (.A(_04712_),
    .B(_04744_),
    .X(_04745_));
 sky130_fd_sc_hd__o211a_1 _10434_ (.A1(\_176_[22] ),
    .A2(_04735_),
    .B1(_04745_),
    .C1(_04740_),
    .X(_00495_));
 sky130_fd_sc_hd__buf_2 _10435_ (.A(_01216_),
    .X(_04746_));
 sky130_fd_sc_hd__or2_1 _10436_ (.A(\_182_[23] ),
    .B(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__o211a_1 _10437_ (.A1(\_179_[23] ),
    .A2(_04721_),
    .B1(_04705_),
    .C1(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__a211o_1 _10438_ (.A1(\_176_[23] ),
    .A2(_04725_),
    .B1(_04748_),
    .C1(_04728_),
    .X(_00496_));
 sky130_fd_sc_hd__or2_1 _10439_ (.A(\_182_[24] ),
    .B(_04746_),
    .X(_04749_));
 sky130_fd_sc_hd__o211a_1 _10440_ (.A1(\_179_[24] ),
    .A2(_04721_),
    .B1(_04705_),
    .C1(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__a211o_1 _10441_ (.A1(\_176_[24] ),
    .A2(_04725_),
    .B1(_04750_),
    .C1(_04728_),
    .X(_00497_));
 sky130_fd_sc_hd__clkbuf_4 _10442_ (.A(_04685_),
    .X(_04751_));
 sky130_fd_sc_hd__or2_1 _10443_ (.A(\_182_[25] ),
    .B(_04746_),
    .X(_04752_));
 sky130_fd_sc_hd__o211a_1 _10444_ (.A1(\_179_[25] ),
    .A2(_04721_),
    .B1(_04751_),
    .C1(_04752_),
    .X(_04753_));
 sky130_fd_sc_hd__a211o_1 _10445_ (.A1(\_176_[25] ),
    .A2(_04725_),
    .B1(_04753_),
    .C1(_04728_),
    .X(_00498_));
 sky130_fd_sc_hd__or2_1 _10446_ (.A(\_182_[26] ),
    .B(_04746_),
    .X(_04754_));
 sky130_fd_sc_hd__o211a_1 _10447_ (.A1(\_179_[26] ),
    .A2(_04721_),
    .B1(_04751_),
    .C1(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__a211o_1 _10448_ (.A1(\_176_[26] ),
    .A2(_04725_),
    .B1(_04755_),
    .C1(_04728_),
    .X(_00499_));
 sky130_fd_sc_hd__or2_1 _10449_ (.A(\_182_[27] ),
    .B(_04746_),
    .X(_04756_));
 sky130_fd_sc_hd__o211a_1 _10450_ (.A1(\_179_[27] ),
    .A2(_04721_),
    .B1(_04751_),
    .C1(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__a211o_1 _10451_ (.A1(\_176_[27] ),
    .A2(_04725_),
    .B1(_04757_),
    .C1(_04728_),
    .X(_00500_));
 sky130_fd_sc_hd__or2_1 _10452_ (.A(\_182_[28] ),
    .B(_04746_),
    .X(_04758_));
 sky130_fd_sc_hd__o211a_1 _10453_ (.A1(\_179_[28] ),
    .A2(_04721_),
    .B1(_04751_),
    .C1(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__a211o_1 _10454_ (.A1(\_176_[28] ),
    .A2(_04725_),
    .B1(_04759_),
    .C1(_04728_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _10455_ (.A0(\_179_[29] ),
    .A1(\_182_[29] ),
    .S(_04743_),
    .X(_04760_));
 sky130_fd_sc_hd__or2_1 _10456_ (.A(_04712_),
    .B(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__o211a_1 _10457_ (.A1(\_176_[29] ),
    .A2(_04735_),
    .B1(_04761_),
    .C1(_04740_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _10458_ (.A0(\_179_[30] ),
    .A1(\_182_[30] ),
    .S(_04743_),
    .X(_04762_));
 sky130_fd_sc_hd__or2_1 _10459_ (.A(_04712_),
    .B(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__o211a_1 _10460_ (.A1(\_176_[30] ),
    .A2(_04735_),
    .B1(_04763_),
    .C1(_04740_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _10461_ (.A0(\_179_[31] ),
    .A1(\_182_[31] ),
    .S(_04743_),
    .X(_04764_));
 sky130_fd_sc_hd__or2_1 _10462_ (.A(_04712_),
    .B(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__o211a_1 _10463_ (.A1(\_176_[31] ),
    .A2(_04735_),
    .B1(_04765_),
    .C1(_04740_),
    .X(_00504_));
 sky130_fd_sc_hd__buf_2 _10464_ (.A(_04681_),
    .X(_04766_));
 sky130_fd_sc_hd__mux2_1 _10465_ (.A0(\_176_[0] ),
    .A1(\_179_[0] ),
    .S(_04743_),
    .X(_04767_));
 sky130_fd_sc_hd__or2_1 _10466_ (.A(_04766_),
    .B(_04767_),
    .X(_04768_));
 sky130_fd_sc_hd__o211a_1 _10467_ (.A1(\_173_[0] ),
    .A2(_04735_),
    .B1(_04768_),
    .C1(_04740_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _10468_ (.A0(\_176_[1] ),
    .A1(\_179_[1] ),
    .S(_04743_),
    .X(_04769_));
 sky130_fd_sc_hd__or2_1 _10469_ (.A(_04766_),
    .B(_04769_),
    .X(_04770_));
 sky130_fd_sc_hd__o211a_1 _10470_ (.A1(\_173_[1] ),
    .A2(_04735_),
    .B1(_04770_),
    .C1(_04740_),
    .X(_00506_));
 sky130_fd_sc_hd__buf_2 _10471_ (.A(_01225_),
    .X(_04771_));
 sky130_fd_sc_hd__or2_1 _10472_ (.A(\_179_[2] ),
    .B(_04746_),
    .X(_04772_));
 sky130_fd_sc_hd__o211a_1 _10473_ (.A1(\_176_[2] ),
    .A2(_04771_),
    .B1(_04751_),
    .C1(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__a211o_1 _10474_ (.A1(\_173_[2] ),
    .A2(_04725_),
    .B1(_04773_),
    .C1(_04728_),
    .X(_00507_));
 sky130_fd_sc_hd__buf_2 _10475_ (.A(_04724_),
    .X(_04774_));
 sky130_fd_sc_hd__or2_1 _10476_ (.A(\_179_[3] ),
    .B(_04746_),
    .X(_04775_));
 sky130_fd_sc_hd__o211a_1 _10477_ (.A1(\_176_[3] ),
    .A2(_04771_),
    .B1(_04751_),
    .C1(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__buf_2 _10478_ (.A(_01418_),
    .X(_04777_));
 sky130_fd_sc_hd__a211o_1 _10479_ (.A1(\_173_[3] ),
    .A2(_04774_),
    .B1(_04776_),
    .C1(_04777_),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _10480_ (.A0(\_176_[4] ),
    .A1(\_179_[4] ),
    .S(_04743_),
    .X(_04778_));
 sky130_fd_sc_hd__or2_1 _10481_ (.A(_04766_),
    .B(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__o211a_1 _10482_ (.A1(\_173_[4] ),
    .A2(_04735_),
    .B1(_04779_),
    .C1(_04740_),
    .X(_00509_));
 sky130_fd_sc_hd__clkbuf_4 _10483_ (.A(_04671_),
    .X(_04780_));
 sky130_fd_sc_hd__mux2_1 _10484_ (.A0(\_176_[5] ),
    .A1(\_179_[5] ),
    .S(_04743_),
    .X(_04781_));
 sky130_fd_sc_hd__or2_1 _10485_ (.A(_04766_),
    .B(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__o211a_1 _10486_ (.A1(\_173_[5] ),
    .A2(_04780_),
    .B1(_04782_),
    .C1(_04740_),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(\_176_[6] ),
    .A1(\_179_[6] ),
    .S(_04743_),
    .X(_04783_));
 sky130_fd_sc_hd__or2_1 _10488_ (.A(_04766_),
    .B(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__clkbuf_4 _10489_ (.A(_01424_),
    .X(_04785_));
 sky130_fd_sc_hd__o211a_1 _10490_ (.A1(\_173_[6] ),
    .A2(_04780_),
    .B1(_04784_),
    .C1(_04785_),
    .X(_00511_));
 sky130_fd_sc_hd__or2_1 _10491_ (.A(\_179_[7] ),
    .B(_04746_),
    .X(_04786_));
 sky130_fd_sc_hd__o211a_1 _10492_ (.A1(\_176_[7] ),
    .A2(_04771_),
    .B1(_04751_),
    .C1(_04786_),
    .X(_04787_));
 sky130_fd_sc_hd__a211o_1 _10493_ (.A1(\_173_[7] ),
    .A2(_04774_),
    .B1(_04787_),
    .C1(_04777_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _10494_ (.A0(\_176_[8] ),
    .A1(\_179_[8] ),
    .S(_04743_),
    .X(_04788_));
 sky130_fd_sc_hd__or2_1 _10495_ (.A(_04766_),
    .B(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__o211a_1 _10496_ (.A1(\_173_[8] ),
    .A2(_04780_),
    .B1(_04789_),
    .C1(_04785_),
    .X(_00513_));
 sky130_fd_sc_hd__buf_4 _10497_ (.A(_01214_),
    .X(_04790_));
 sky130_fd_sc_hd__mux2_1 _10498_ (.A0(\_176_[9] ),
    .A1(\_179_[9] ),
    .S(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__or2_1 _10499_ (.A(_04766_),
    .B(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__o211a_1 _10500_ (.A1(\_173_[9] ),
    .A2(_04780_),
    .B1(_04792_),
    .C1(_04785_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _10501_ (.A0(\_176_[10] ),
    .A1(\_179_[10] ),
    .S(_04790_),
    .X(_04793_));
 sky130_fd_sc_hd__or2_1 _10502_ (.A(_04766_),
    .B(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__o211a_1 _10503_ (.A1(\_173_[10] ),
    .A2(_04780_),
    .B1(_04794_),
    .C1(_04785_),
    .X(_00515_));
 sky130_fd_sc_hd__or2_1 _10504_ (.A(\_179_[11] ),
    .B(_04746_),
    .X(_04795_));
 sky130_fd_sc_hd__o211a_1 _10505_ (.A1(\_176_[11] ),
    .A2(_04771_),
    .B1(_04751_),
    .C1(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__a211o_1 _10506_ (.A1(\_173_[11] ),
    .A2(_04774_),
    .B1(_04796_),
    .C1(_04777_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _10507_ (.A0(\_176_[12] ),
    .A1(\_179_[12] ),
    .S(_04790_),
    .X(_04797_));
 sky130_fd_sc_hd__or2_1 _10508_ (.A(_04766_),
    .B(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__o211a_1 _10509_ (.A1(\_173_[12] ),
    .A2(_04780_),
    .B1(_04798_),
    .C1(_04785_),
    .X(_00517_));
 sky130_fd_sc_hd__clkbuf_2 _10510_ (.A(_01216_),
    .X(_04799_));
 sky130_fd_sc_hd__or2_1 _10511_ (.A(\_179_[13] ),
    .B(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__o211a_1 _10512_ (.A1(\_176_[13] ),
    .A2(_04771_),
    .B1(_04751_),
    .C1(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__a211o_1 _10513_ (.A1(\_173_[13] ),
    .A2(_04774_),
    .B1(_04801_),
    .C1(_04777_),
    .X(_00518_));
 sky130_fd_sc_hd__or2_1 _10514_ (.A(\_179_[14] ),
    .B(_04799_),
    .X(_04802_));
 sky130_fd_sc_hd__o211a_1 _10515_ (.A1(\_176_[14] ),
    .A2(_04771_),
    .B1(_04751_),
    .C1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__a211o_1 _10516_ (.A1(\_173_[14] ),
    .A2(_04774_),
    .B1(_04803_),
    .C1(_04777_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(\_176_[15] ),
    .A1(\_179_[15] ),
    .S(_04790_),
    .X(_04804_));
 sky130_fd_sc_hd__or2_1 _10518_ (.A(_04766_),
    .B(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__o211a_1 _10519_ (.A1(\_173_[15] ),
    .A2(_04780_),
    .B1(_04805_),
    .C1(_04785_),
    .X(_00520_));
 sky130_fd_sc_hd__buf_2 _10520_ (.A(_04685_),
    .X(_04806_));
 sky130_fd_sc_hd__or2_1 _10521_ (.A(\_179_[16] ),
    .B(_04799_),
    .X(_04807_));
 sky130_fd_sc_hd__o211a_1 _10522_ (.A1(\_176_[16] ),
    .A2(_04771_),
    .B1(_04806_),
    .C1(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__a211o_1 _10523_ (.A1(\_173_[16] ),
    .A2(_04774_),
    .B1(_04808_),
    .C1(_04777_),
    .X(_00521_));
 sky130_fd_sc_hd__buf_2 _10524_ (.A(_04681_),
    .X(_04809_));
 sky130_fd_sc_hd__mux2_1 _10525_ (.A0(\_176_[17] ),
    .A1(\_179_[17] ),
    .S(_04790_),
    .X(_04810_));
 sky130_fd_sc_hd__or2_1 _10526_ (.A(_04809_),
    .B(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__o211a_1 _10527_ (.A1(\_173_[17] ),
    .A2(_04780_),
    .B1(_04811_),
    .C1(_04785_),
    .X(_00522_));
 sky130_fd_sc_hd__or2_1 _10528_ (.A(\_179_[18] ),
    .B(_04799_),
    .X(_04812_));
 sky130_fd_sc_hd__o211a_1 _10529_ (.A1(\_176_[18] ),
    .A2(_04771_),
    .B1(_04806_),
    .C1(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__a211o_1 _10530_ (.A1(\_173_[18] ),
    .A2(_04774_),
    .B1(_04813_),
    .C1(_04777_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _10531_ (.A0(\_176_[19] ),
    .A1(\_179_[19] ),
    .S(_04790_),
    .X(_04814_));
 sky130_fd_sc_hd__or2_1 _10532_ (.A(_04809_),
    .B(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__o211a_1 _10533_ (.A1(\_173_[19] ),
    .A2(_04780_),
    .B1(_04815_),
    .C1(_04785_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _10534_ (.A0(\_176_[20] ),
    .A1(\_179_[20] ),
    .S(_04790_),
    .X(_04816_));
 sky130_fd_sc_hd__or2_1 _10535_ (.A(_04809_),
    .B(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__o211a_1 _10536_ (.A1(\_173_[20] ),
    .A2(_04780_),
    .B1(_04817_),
    .C1(_04785_),
    .X(_00525_));
 sky130_fd_sc_hd__clkbuf_4 _10537_ (.A(_04671_),
    .X(_04818_));
 sky130_fd_sc_hd__mux2_1 _10538_ (.A0(\_176_[21] ),
    .A1(\_179_[21] ),
    .S(_04790_),
    .X(_04819_));
 sky130_fd_sc_hd__or2_1 _10539_ (.A(_04809_),
    .B(_04819_),
    .X(_04820_));
 sky130_fd_sc_hd__o211a_1 _10540_ (.A1(\_173_[21] ),
    .A2(_04818_),
    .B1(_04820_),
    .C1(_04785_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _10541_ (.A0(\_176_[22] ),
    .A1(\_179_[22] ),
    .S(_04790_),
    .X(_04821_));
 sky130_fd_sc_hd__or2_1 _10542_ (.A(_04809_),
    .B(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__clkbuf_4 _10543_ (.A(_01424_),
    .X(_04823_));
 sky130_fd_sc_hd__o211a_1 _10544_ (.A1(\_173_[22] ),
    .A2(_04818_),
    .B1(_04822_),
    .C1(_04823_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _10545_ (.A0(\_176_[23] ),
    .A1(\_179_[23] ),
    .S(_04790_),
    .X(_04824_));
 sky130_fd_sc_hd__or2_1 _10546_ (.A(_04809_),
    .B(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__o211a_1 _10547_ (.A1(\_173_[23] ),
    .A2(_04818_),
    .B1(_04825_),
    .C1(_04823_),
    .X(_00528_));
 sky130_fd_sc_hd__or2_1 _10548_ (.A(\_179_[24] ),
    .B(_04799_),
    .X(_04826_));
 sky130_fd_sc_hd__o211a_1 _10549_ (.A1(\_176_[24] ),
    .A2(_04771_),
    .B1(_04806_),
    .C1(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__a211o_1 _10550_ (.A1(\_173_[24] ),
    .A2(_04774_),
    .B1(_04827_),
    .C1(_04777_),
    .X(_00529_));
 sky130_fd_sc_hd__or2_1 _10551_ (.A(\_179_[25] ),
    .B(_04799_),
    .X(_04828_));
 sky130_fd_sc_hd__o211a_1 _10552_ (.A1(\_176_[25] ),
    .A2(_04771_),
    .B1(_04806_),
    .C1(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__a211o_1 _10553_ (.A1(\_173_[25] ),
    .A2(_04774_),
    .B1(_04829_),
    .C1(_04777_),
    .X(_00530_));
 sky130_fd_sc_hd__clkbuf_4 _10554_ (.A(_01213_),
    .X(_04830_));
 sky130_fd_sc_hd__mux2_1 _10555_ (.A0(\_176_[26] ),
    .A1(\_179_[26] ),
    .S(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__or2_1 _10556_ (.A(_04809_),
    .B(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__o211a_1 _10557_ (.A1(\_173_[26] ),
    .A2(_04818_),
    .B1(_04832_),
    .C1(_04823_),
    .X(_00531_));
 sky130_fd_sc_hd__clkbuf_4 _10558_ (.A(_01225_),
    .X(_04833_));
 sky130_fd_sc_hd__or2_1 _10559_ (.A(\_179_[27] ),
    .B(_04799_),
    .X(_04834_));
 sky130_fd_sc_hd__o211a_1 _10560_ (.A1(\_176_[27] ),
    .A2(_04833_),
    .B1(_04806_),
    .C1(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__a211o_1 _10561_ (.A1(\_173_[27] ),
    .A2(_04774_),
    .B1(_04835_),
    .C1(_04777_),
    .X(_00532_));
 sky130_fd_sc_hd__clkbuf_4 _10562_ (.A(_04682_),
    .X(_04836_));
 sky130_fd_sc_hd__or2_1 _10563_ (.A(\_179_[28] ),
    .B(_04799_),
    .X(_04837_));
 sky130_fd_sc_hd__o211a_1 _10564_ (.A1(\_176_[28] ),
    .A2(_04833_),
    .B1(_04806_),
    .C1(_04837_),
    .X(_04838_));
 sky130_fd_sc_hd__clkbuf_4 _10565_ (.A(_01418_),
    .X(_04839_));
 sky130_fd_sc_hd__a211o_1 _10566_ (.A1(\_173_[28] ),
    .A2(_04836_),
    .B1(_04838_),
    .C1(_04839_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _10567_ (.A0(\_176_[29] ),
    .A1(\_179_[29] ),
    .S(_04830_),
    .X(_04840_));
 sky130_fd_sc_hd__or2_1 _10568_ (.A(_04809_),
    .B(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__o211a_1 _10569_ (.A1(\_173_[29] ),
    .A2(_04818_),
    .B1(_04841_),
    .C1(_04823_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(\_176_[30] ),
    .A1(\_179_[30] ),
    .S(_04830_),
    .X(_04842_));
 sky130_fd_sc_hd__or2_1 _10571_ (.A(_04809_),
    .B(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__o211a_1 _10572_ (.A1(\_173_[30] ),
    .A2(_04818_),
    .B1(_04843_),
    .C1(_04823_),
    .X(_00535_));
 sky130_fd_sc_hd__or2_1 _10573_ (.A(\_179_[31] ),
    .B(_04799_),
    .X(_04844_));
 sky130_fd_sc_hd__o211a_1 _10574_ (.A1(\_176_[31] ),
    .A2(_04833_),
    .B1(_04806_),
    .C1(_04844_),
    .X(_04845_));
 sky130_fd_sc_hd__a211o_1 _10575_ (.A1(\_173_[31] ),
    .A2(_04836_),
    .B1(_04845_),
    .C1(_04839_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _10576_ (.A0(\_173_[0] ),
    .A1(\_176_[0] ),
    .S(_01226_),
    .X(_04846_));
 sky130_fd_sc_hd__a31o_1 _10577_ (.A1(_01711_),
    .A2(_01712_),
    .A3(_04724_),
    .B1(_01710_),
    .X(_04847_));
 sky130_fd_sc_hd__a21o_1 _10578_ (.A1(_04691_),
    .A2(_04846_),
    .B1(_04847_),
    .X(_00537_));
 sky130_fd_sc_hd__buf_4 _10579_ (.A(_04637_),
    .X(_04848_));
 sky130_fd_sc_hd__clkbuf_4 _10580_ (.A(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__a221o_1 _10581_ (.A1(\_176_[1] ),
    .A2(net68),
    .B1(_01741_),
    .B2(_04682_),
    .C1(_02711_),
    .X(_04850_));
 sky130_fd_sc_hd__a21o_1 _10582_ (.A1(\_173_[1] ),
    .A2(_04849_),
    .B1(_04850_),
    .X(_00538_));
 sky130_fd_sc_hd__a221o_1 _10583_ (.A1(\_176_[2] ),
    .A2(net68),
    .B1(_01751_),
    .B2(_04682_),
    .C1(_02711_),
    .X(_04851_));
 sky130_fd_sc_hd__a21o_1 _10584_ (.A1(\_173_[2] ),
    .A2(_04849_),
    .B1(_04851_),
    .X(_00539_));
 sky130_fd_sc_hd__a221o_1 _10585_ (.A1(\_176_[3] ),
    .A2(net68),
    .B1(_01777_),
    .B2(_04692_),
    .C1(_02711_),
    .X(_04852_));
 sky130_fd_sc_hd__a21o_1 _10586_ (.A1(\_173_[3] ),
    .A2(_04849_),
    .B1(_04852_),
    .X(_00540_));
 sky130_fd_sc_hd__buf_4 _10587_ (.A(_04686_),
    .X(_04853_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(\_173_[4] ),
    .A1(\_176_[4] ),
    .S(_01226_),
    .X(_04854_));
 sky130_fd_sc_hd__buf_4 _10589_ (.A(_04630_),
    .X(_04855_));
 sky130_fd_sc_hd__nor2_1 _10590_ (.A(_01824_),
    .B(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__a211o_1 _10591_ (.A1(_04853_),
    .A2(_04854_),
    .B1(_04856_),
    .C1(_04839_),
    .X(_00541_));
 sky130_fd_sc_hd__a221o_1 _10592_ (.A1(\_176_[5] ),
    .A2(net68),
    .B1(_01833_),
    .B2(_04692_),
    .C1(_02711_),
    .X(_04857_));
 sky130_fd_sc_hd__a21o_1 _10593_ (.A1(\_173_[5] ),
    .A2(_04849_),
    .B1(_04857_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _10594_ (.A0(\_173_[6] ),
    .A1(\_176_[6] ),
    .S(_01226_),
    .X(_04858_));
 sky130_fd_sc_hd__nor2_1 _10595_ (.A(_01863_),
    .B(_04631_),
    .Y(_04859_));
 sky130_fd_sc_hd__a211o_1 _10596_ (.A1(_04853_),
    .A2(_04858_),
    .B1(_04859_),
    .C1(_04839_),
    .X(_00543_));
 sky130_fd_sc_hd__o221a_1 _10597_ (.A1(\_176_[7] ),
    .A2(_04678_),
    .B1(_01892_),
    .B2(_04686_),
    .C1(_04648_),
    .X(_04860_));
 sky130_fd_sc_hd__o21a_1 _10598_ (.A1(\_173_[7] ),
    .A2(_04629_),
    .B1(_04860_),
    .X(_00544_));
 sky130_fd_sc_hd__buf_6 _10599_ (.A(_04724_),
    .X(_04861_));
 sky130_fd_sc_hd__mux2_1 _10600_ (.A0(\_173_[8] ),
    .A1(\_176_[8] ),
    .S(_01226_),
    .X(_04862_));
 sky130_fd_sc_hd__nand2_1 _10601_ (.A(_01922_),
    .B(_04724_),
    .Y(_04863_));
 sky130_fd_sc_hd__o211a_1 _10602_ (.A1(_04861_),
    .A2(_04862_),
    .B1(_04863_),
    .C1(_04823_),
    .X(_00545_));
 sky130_fd_sc_hd__inv_2 _10603_ (.A(\_176_[9] ),
    .Y(_04864_));
 sky130_fd_sc_hd__buf_4 _10604_ (.A(_04625_),
    .X(_04865_));
 sky130_fd_sc_hd__o221a_1 _10605_ (.A1(_04864_),
    .A2(_04678_),
    .B1(_01971_),
    .B2(_04865_),
    .C1(_02833_),
    .X(_04866_));
 sky130_fd_sc_hd__a21bo_1 _10606_ (.A1(\_173_[9] ),
    .A2(_04849_),
    .B1_N(_04866_),
    .X(_00546_));
 sky130_fd_sc_hd__buf_4 _10607_ (.A(_01212_),
    .X(_04867_));
 sky130_fd_sc_hd__or2_1 _10608_ (.A(\_176_[10] ),
    .B(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__mux2_1 _10609_ (.A0(_02001_),
    .A1(_04868_),
    .S(_04865_),
    .X(_04869_));
 sky130_fd_sc_hd__o211a_1 _10610_ (.A1(\_173_[10] ),
    .A2(_04663_),
    .B1(_04869_),
    .C1(_04823_),
    .X(_00547_));
 sky130_fd_sc_hd__or2_1 _10611_ (.A(\_176_[11] ),
    .B(_04867_),
    .X(_04870_));
 sky130_fd_sc_hd__mux2_1 _10612_ (.A0(_02028_),
    .A1(_04870_),
    .S(_04630_),
    .X(_04871_));
 sky130_fd_sc_hd__o211a_1 _10613_ (.A1(\_173_[11] ),
    .A2(_04663_),
    .B1(_04871_),
    .C1(_04823_),
    .X(_00548_));
 sky130_fd_sc_hd__buf_4 _10614_ (.A(_04636_),
    .X(_04872_));
 sky130_fd_sc_hd__nand2_1 _10615_ (.A(_02058_),
    .B(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__o211a_1 _10616_ (.A1(\_176_[12] ),
    .A2(_04872_),
    .B1(_04633_),
    .C1(_04873_),
    .X(_04874_));
 sky130_fd_sc_hd__a211o_1 _10617_ (.A1(\_173_[12] ),
    .A2(_04849_),
    .B1(_04874_),
    .C1(_04839_),
    .X(_00549_));
 sky130_fd_sc_hd__o221a_1 _10618_ (.A1(\_176_[13] ),
    .A2(_04678_),
    .B1(_04627_),
    .B2(\_173_[13] ),
    .C1(_02833_),
    .X(_04875_));
 sky130_fd_sc_hd__a21boi_1 _10619_ (.A1(_02085_),
    .A2(_04861_),
    .B1_N(_04875_),
    .Y(_00550_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(\_173_[14] ),
    .A1(\_176_[14] ),
    .S(_01215_),
    .X(_04876_));
 sky130_fd_sc_hd__nor2_1 _10621_ (.A(_02111_),
    .B(_04631_),
    .Y(_04877_));
 sky130_fd_sc_hd__a211o_1 _10622_ (.A1(_04853_),
    .A2(_04876_),
    .B1(_04877_),
    .C1(_04839_),
    .X(_00551_));
 sky130_fd_sc_hd__o221a_1 _10623_ (.A1(\_176_[15] ),
    .A2(_04678_),
    .B1(_04627_),
    .B2(\_173_[15] ),
    .C1(_02833_),
    .X(_04878_));
 sky130_fd_sc_hd__a21boi_1 _10624_ (.A1(_02139_),
    .A2(_04861_),
    .B1_N(_04878_),
    .Y(_00552_));
 sky130_fd_sc_hd__mux2_1 _10625_ (.A0(\_173_[16] ),
    .A1(\_176_[16] ),
    .S(_04830_),
    .X(_04879_));
 sky130_fd_sc_hd__or2_1 _10626_ (.A(_04809_),
    .B(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__o211a_1 _10627_ (.A1(_02175_),
    .A2(_04818_),
    .B1(_04880_),
    .C1(_04823_),
    .X(_00553_));
 sky130_fd_sc_hd__a21o_1 _10628_ (.A1(\_176_[17] ),
    .A2(_04684_),
    .B1(_01417_),
    .X(_04881_));
 sky130_fd_sc_hd__a221o_1 _10629_ (.A1(_02181_),
    .A2(_04724_),
    .B1(_04848_),
    .B2(\_173_[17] ),
    .C1(_04881_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(\_173_[18] ),
    .A1(\_176_[18] ),
    .S(_01215_),
    .X(_04882_));
 sky130_fd_sc_hd__nor2_1 _10631_ (.A(_02230_),
    .B(_04631_),
    .Y(_04883_));
 sky130_fd_sc_hd__a211o_1 _10632_ (.A1(_04855_),
    .A2(_04882_),
    .B1(_04883_),
    .C1(_04839_),
    .X(_00555_));
 sky130_fd_sc_hd__or2_1 _10633_ (.A(_02237_),
    .B(_04685_),
    .X(_04884_));
 sky130_fd_sc_hd__o211a_1 _10634_ (.A1(\_176_[19] ),
    .A2(_04872_),
    .B1(_04633_),
    .C1(_04884_),
    .X(_04885_));
 sky130_fd_sc_hd__a211o_1 _10635_ (.A1(\_173_[19] ),
    .A2(_04848_),
    .B1(_04885_),
    .C1(_04839_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _10636_ (.A0(\_173_[20] ),
    .A1(\_176_[20] ),
    .S(_01226_),
    .X(_04886_));
 sky130_fd_sc_hd__nand2_1 _10637_ (.A(_02293_),
    .B(_04724_),
    .Y(_04887_));
 sky130_fd_sc_hd__o211a_1 _10638_ (.A1(_04861_),
    .A2(_04886_),
    .B1(_04887_),
    .C1(_04823_),
    .X(_00557_));
 sky130_fd_sc_hd__clkbuf_2 _10639_ (.A(_04681_),
    .X(_04888_));
 sky130_fd_sc_hd__mux2_1 _10640_ (.A0(\_173_[21] ),
    .A1(\_176_[21] ),
    .S(_04830_),
    .X(_04889_));
 sky130_fd_sc_hd__or2_1 _10641_ (.A(_04888_),
    .B(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__clkbuf_4 _10642_ (.A(_01424_),
    .X(_04891_));
 sky130_fd_sc_hd__o211a_1 _10643_ (.A1(_02300_),
    .A2(_04818_),
    .B1(_04890_),
    .C1(_04891_),
    .X(_00558_));
 sky130_fd_sc_hd__or2_1 _10644_ (.A(\_176_[22] ),
    .B(_04867_),
    .X(_04892_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(_02353_),
    .A1(_04892_),
    .S(_04630_),
    .X(_04893_));
 sky130_fd_sc_hd__o211a_1 _10646_ (.A1(\_173_[22] ),
    .A2(_04663_),
    .B1(_04893_),
    .C1(_04891_),
    .X(_00559_));
 sky130_fd_sc_hd__or2_1 _10647_ (.A(\_176_[23] ),
    .B(_01216_),
    .X(_04894_));
 sky130_fd_sc_hd__mux2_1 _10648_ (.A0(_02359_),
    .A1(_04894_),
    .S(_04630_),
    .X(_04895_));
 sky130_fd_sc_hd__o211a_1 _10649_ (.A1(\_173_[23] ),
    .A2(_04663_),
    .B1(_04895_),
    .C1(_04891_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(\_173_[24] ),
    .A1(\_176_[24] ),
    .S(_01215_),
    .X(_04896_));
 sky130_fd_sc_hd__nor2_1 _10651_ (.A(_02416_),
    .B(_04631_),
    .Y(_04897_));
 sky130_fd_sc_hd__a211o_1 _10652_ (.A1(_04855_),
    .A2(_04896_),
    .B1(_04897_),
    .C1(_04839_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _10653_ (.A0(\_173_[25] ),
    .A1(\_176_[25] ),
    .S(_01226_),
    .X(_04898_));
 sky130_fd_sc_hd__nand2_1 _10654_ (.A(_02445_),
    .B(_04724_),
    .Y(_04899_));
 sky130_fd_sc_hd__o211a_1 _10655_ (.A1(_04861_),
    .A2(_04898_),
    .B1(_04899_),
    .C1(_04891_),
    .X(_00562_));
 sky130_fd_sc_hd__o221a_1 _10656_ (.A1(\_176_[26] ),
    .A2(_04678_),
    .B1(_04627_),
    .B2(\_173_[26] ),
    .C1(_02833_),
    .X(_04900_));
 sky130_fd_sc_hd__a21boi_1 _10657_ (.A1(_02476_),
    .A2(_04861_),
    .B1_N(_04900_),
    .Y(_00563_));
 sky130_fd_sc_hd__o221a_1 _10658_ (.A1(\_176_[27] ),
    .A2(_04678_),
    .B1(_04633_),
    .B2(\_173_[27] ),
    .C1(_04648_),
    .X(_04901_));
 sky130_fd_sc_hd__o21a_1 _10659_ (.A1(_02483_),
    .A2(_04691_),
    .B1(_04901_),
    .X(_00564_));
 sky130_fd_sc_hd__nand2_1 _10660_ (.A(_02535_),
    .B(_04872_),
    .Y(_04902_));
 sky130_fd_sc_hd__o211a_1 _10661_ (.A1(\_176_[28] ),
    .A2(_04872_),
    .B1(_04633_),
    .C1(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__a211o_1 _10662_ (.A1(\_173_[28] ),
    .A2(_04848_),
    .B1(_04903_),
    .C1(_04839_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _10663_ (.A0(\_173_[29] ),
    .A1(\_176_[29] ),
    .S(_01226_),
    .X(_04904_));
 sky130_fd_sc_hd__nand2_1 _10664_ (.A(_02561_),
    .B(_04724_),
    .Y(_04905_));
 sky130_fd_sc_hd__o211a_1 _10665_ (.A1(_04683_),
    .A2(_04904_),
    .B1(_04905_),
    .C1(_04891_),
    .X(_00566_));
 sky130_fd_sc_hd__a221o_1 _10666_ (.A1(\_176_[30] ),
    .A2(net68),
    .B1(_04638_),
    .B2(\_173_[30] ),
    .C1(_02711_),
    .X(_04906_));
 sky130_fd_sc_hd__a21o_1 _10667_ (.A1(_02570_),
    .A2(_04861_),
    .B1(_04906_),
    .X(_00567_));
 sky130_fd_sc_hd__nand2_1 _10668_ (.A(\_173_[31] ),
    .B(_04848_),
    .Y(_04907_));
 sky130_fd_sc_hd__nor2_1 _10669_ (.A(\_176_[31] ),
    .B(_04681_),
    .Y(_04908_));
 sky130_fd_sc_hd__a211o_1 _10670_ (.A1(_02606_),
    .A2(_04872_),
    .B1(_04637_),
    .C1(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__a21oi_1 _10671_ (.A1(_04907_),
    .A2(_04909_),
    .B1(_03866_),
    .Y(_00568_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(\_170_[0] ),
    .A1(\_173_[0] ),
    .S(_04830_),
    .X(_04910_));
 sky130_fd_sc_hd__or2_1 _10673_ (.A(_04888_),
    .B(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__o211a_1 _10674_ (.A1(\_167_[0] ),
    .A2(_04818_),
    .B1(_04911_),
    .C1(_04891_),
    .X(_00569_));
 sky130_fd_sc_hd__or2_1 _10675_ (.A(\_173_[1] ),
    .B(_04799_),
    .X(_04912_));
 sky130_fd_sc_hd__o211a_1 _10676_ (.A1(\_170_[1] ),
    .A2(_04833_),
    .B1(_04806_),
    .C1(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__buf_2 _10677_ (.A(_01418_),
    .X(_04914_));
 sky130_fd_sc_hd__a211o_1 _10678_ (.A1(\_167_[1] ),
    .A2(_04836_),
    .B1(_04913_),
    .C1(_04914_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _10679_ (.A0(\_170_[2] ),
    .A1(\_173_[2] ),
    .S(_04830_),
    .X(_04915_));
 sky130_fd_sc_hd__or2_1 _10680_ (.A(_04888_),
    .B(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__o211a_1 _10681_ (.A1(\_167_[2] ),
    .A2(_04818_),
    .B1(_04916_),
    .C1(_04891_),
    .X(_00571_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10682_ (.A(_01216_),
    .X(_04917_));
 sky130_fd_sc_hd__or2_1 _10683_ (.A(\_173_[3] ),
    .B(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__o211a_1 _10684_ (.A1(\_170_[3] ),
    .A2(_04833_),
    .B1(_04806_),
    .C1(_04918_),
    .X(_04919_));
 sky130_fd_sc_hd__a211o_1 _10685_ (.A1(\_167_[3] ),
    .A2(_04836_),
    .B1(_04919_),
    .C1(_04914_),
    .X(_00572_));
 sky130_fd_sc_hd__or2_1 _10686_ (.A(\_173_[4] ),
    .B(_04917_),
    .X(_04920_));
 sky130_fd_sc_hd__o211a_1 _10687_ (.A1(\_170_[4] ),
    .A2(_04833_),
    .B1(_04806_),
    .C1(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__a211o_1 _10688_ (.A1(\_167_[4] ),
    .A2(_04836_),
    .B1(_04921_),
    .C1(_04914_),
    .X(_00573_));
 sky130_fd_sc_hd__buf_2 _10689_ (.A(_04685_),
    .X(_04922_));
 sky130_fd_sc_hd__or2_1 _10690_ (.A(\_173_[5] ),
    .B(_04917_),
    .X(_04923_));
 sky130_fd_sc_hd__o211a_1 _10691_ (.A1(\_170_[5] ),
    .A2(_04833_),
    .B1(_04922_),
    .C1(_04923_),
    .X(_04924_));
 sky130_fd_sc_hd__a211o_1 _10692_ (.A1(\_167_[5] ),
    .A2(_04836_),
    .B1(_04924_),
    .C1(_04914_),
    .X(_00574_));
 sky130_fd_sc_hd__clkbuf_4 _10693_ (.A(_04671_),
    .X(_04925_));
 sky130_fd_sc_hd__mux2_1 _10694_ (.A0(\_170_[6] ),
    .A1(\_173_[6] ),
    .S(_04830_),
    .X(_04926_));
 sky130_fd_sc_hd__or2_1 _10695_ (.A(_04888_),
    .B(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__o211a_1 _10696_ (.A1(\_167_[6] ),
    .A2(_04925_),
    .B1(_04927_),
    .C1(_04891_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _10697_ (.A0(\_170_[7] ),
    .A1(\_173_[7] ),
    .S(_04830_),
    .X(_04928_));
 sky130_fd_sc_hd__or2_1 _10698_ (.A(_04888_),
    .B(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__o211a_1 _10699_ (.A1(\_167_[7] ),
    .A2(_04925_),
    .B1(_04929_),
    .C1(_04891_),
    .X(_00576_));
 sky130_fd_sc_hd__or2_1 _10700_ (.A(\_173_[8] ),
    .B(_04917_),
    .X(_04930_));
 sky130_fd_sc_hd__o211a_1 _10701_ (.A1(\_170_[8] ),
    .A2(_04833_),
    .B1(_04922_),
    .C1(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__a211o_1 _10702_ (.A1(\_167_[8] ),
    .A2(_04836_),
    .B1(_04931_),
    .C1(_04914_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _10703_ (.A0(\_170_[9] ),
    .A1(\_173_[9] ),
    .S(_04830_),
    .X(_04932_));
 sky130_fd_sc_hd__or2_1 _10704_ (.A(_04888_),
    .B(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__o211a_1 _10705_ (.A1(\_167_[9] ),
    .A2(_04925_),
    .B1(_04933_),
    .C1(_04891_),
    .X(_00578_));
 sky130_fd_sc_hd__or2_1 _10706_ (.A(\_173_[10] ),
    .B(_04917_),
    .X(_04934_));
 sky130_fd_sc_hd__o211a_1 _10707_ (.A1(\_170_[10] ),
    .A2(_04833_),
    .B1(_04922_),
    .C1(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__a211o_1 _10708_ (.A1(\_167_[10] ),
    .A2(_04836_),
    .B1(_04935_),
    .C1(_04914_),
    .X(_00579_));
 sky130_fd_sc_hd__clkbuf_4 _10709_ (.A(_01213_),
    .X(_04936_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(\_170_[11] ),
    .A1(\_173_[11] ),
    .S(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__or2_1 _10711_ (.A(_04888_),
    .B(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__buf_2 _10712_ (.A(_01424_),
    .X(_04939_));
 sky130_fd_sc_hd__o211a_1 _10713_ (.A1(\_167_[11] ),
    .A2(_04925_),
    .B1(_04938_),
    .C1(_04939_),
    .X(_00580_));
 sky130_fd_sc_hd__or2_1 _10714_ (.A(\_173_[12] ),
    .B(_04917_),
    .X(_04940_));
 sky130_fd_sc_hd__o211a_1 _10715_ (.A1(\_170_[12] ),
    .A2(_04833_),
    .B1(_04922_),
    .C1(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__a211o_1 _10716_ (.A1(\_167_[12] ),
    .A2(_04836_),
    .B1(_04941_),
    .C1(_04914_),
    .X(_00581_));
 sky130_fd_sc_hd__buf_2 _10717_ (.A(_01225_),
    .X(_04942_));
 sky130_fd_sc_hd__or2_1 _10718_ (.A(\_173_[13] ),
    .B(_04917_),
    .X(_04943_));
 sky130_fd_sc_hd__o211a_1 _10719_ (.A1(\_170_[13] ),
    .A2(_04942_),
    .B1(_04922_),
    .C1(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__a211o_1 _10720_ (.A1(\_167_[13] ),
    .A2(_04836_),
    .B1(_04944_),
    .C1(_04914_),
    .X(_00582_));
 sky130_fd_sc_hd__buf_2 _10721_ (.A(_04682_),
    .X(_04945_));
 sky130_fd_sc_hd__or2_1 _10722_ (.A(\_173_[14] ),
    .B(_04917_),
    .X(_04946_));
 sky130_fd_sc_hd__o211a_1 _10723_ (.A1(\_170_[14] ),
    .A2(_04942_),
    .B1(_04922_),
    .C1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__a211o_1 _10724_ (.A1(\_167_[14] ),
    .A2(_04945_),
    .B1(_04947_),
    .C1(_04914_),
    .X(_00583_));
 sky130_fd_sc_hd__or2_1 _10725_ (.A(\_173_[15] ),
    .B(_04917_),
    .X(_04948_));
 sky130_fd_sc_hd__o211a_1 _10726_ (.A1(\_170_[15] ),
    .A2(_04942_),
    .B1(_04922_),
    .C1(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__a211o_1 _10727_ (.A1(\_167_[15] ),
    .A2(_04945_),
    .B1(_04949_),
    .C1(_04914_),
    .X(_00584_));
 sky130_fd_sc_hd__or2_1 _10728_ (.A(\_173_[16] ),
    .B(_04917_),
    .X(_04950_));
 sky130_fd_sc_hd__o211a_1 _10729_ (.A1(\_170_[16] ),
    .A2(_04942_),
    .B1(_04922_),
    .C1(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__clkbuf_4 _10730_ (.A(_01418_),
    .X(_04952_));
 sky130_fd_sc_hd__a211o_1 _10731_ (.A1(\_167_[16] ),
    .A2(_04945_),
    .B1(_04951_),
    .C1(_04952_),
    .X(_00585_));
 sky130_fd_sc_hd__clkbuf_2 _10732_ (.A(_01216_),
    .X(_04953_));
 sky130_fd_sc_hd__or2_1 _10733_ (.A(\_173_[17] ),
    .B(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__o211a_1 _10734_ (.A1(\_170_[17] ),
    .A2(_04942_),
    .B1(_04922_),
    .C1(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__a211o_1 _10735_ (.A1(\_167_[17] ),
    .A2(_04945_),
    .B1(_04955_),
    .C1(_04952_),
    .X(_00586_));
 sky130_fd_sc_hd__or2_1 _10736_ (.A(\_173_[18] ),
    .B(_04953_),
    .X(_04956_));
 sky130_fd_sc_hd__o211a_1 _10737_ (.A1(\_170_[18] ),
    .A2(_04942_),
    .B1(_04922_),
    .C1(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__a211o_1 _10738_ (.A1(\_167_[18] ),
    .A2(_04945_),
    .B1(_04957_),
    .C1(_04952_),
    .X(_00587_));
 sky130_fd_sc_hd__clkbuf_4 _10739_ (.A(_04685_),
    .X(_04958_));
 sky130_fd_sc_hd__or2_1 _10740_ (.A(\_173_[19] ),
    .B(_04953_),
    .X(_04959_));
 sky130_fd_sc_hd__o211a_1 _10741_ (.A1(\_170_[19] ),
    .A2(_04942_),
    .B1(_04958_),
    .C1(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__a211o_1 _10742_ (.A1(\_167_[19] ),
    .A2(_04945_),
    .B1(_04960_),
    .C1(_04952_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\_170_[20] ),
    .A1(\_173_[20] ),
    .S(_04936_),
    .X(_04961_));
 sky130_fd_sc_hd__or2_1 _10744_ (.A(_04888_),
    .B(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__o211a_1 _10745_ (.A1(\_167_[20] ),
    .A2(_04925_),
    .B1(_04962_),
    .C1(_04939_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(\_170_[21] ),
    .A1(\_173_[21] ),
    .S(_04936_),
    .X(_04963_));
 sky130_fd_sc_hd__or2_1 _10747_ (.A(_04888_),
    .B(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__o211a_1 _10748_ (.A1(\_167_[21] ),
    .A2(_04925_),
    .B1(_04964_),
    .C1(_04939_),
    .X(_00590_));
 sky130_fd_sc_hd__or2_1 _10749_ (.A(\_173_[22] ),
    .B(_04953_),
    .X(_04965_));
 sky130_fd_sc_hd__o211a_1 _10750_ (.A1(\_170_[22] ),
    .A2(_04942_),
    .B1(_04958_),
    .C1(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__a211o_1 _10751_ (.A1(\_167_[22] ),
    .A2(_04945_),
    .B1(_04966_),
    .C1(_04952_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(\_170_[23] ),
    .A1(\_173_[23] ),
    .S(_04936_),
    .X(_04967_));
 sky130_fd_sc_hd__or2_1 _10753_ (.A(_04888_),
    .B(_04967_),
    .X(_04968_));
 sky130_fd_sc_hd__o211a_1 _10754_ (.A1(\_167_[23] ),
    .A2(_04925_),
    .B1(_04968_),
    .C1(_04939_),
    .X(_00592_));
 sky130_fd_sc_hd__or2_1 _10755_ (.A(\_173_[24] ),
    .B(_04953_),
    .X(_04969_));
 sky130_fd_sc_hd__o211a_1 _10756_ (.A1(\_170_[24] ),
    .A2(_04942_),
    .B1(_04958_),
    .C1(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__a211o_1 _10757_ (.A1(\_167_[24] ),
    .A2(_04945_),
    .B1(_04970_),
    .C1(_04952_),
    .X(_00593_));
 sky130_fd_sc_hd__clkbuf_2 _10758_ (.A(_04636_),
    .X(_04971_));
 sky130_fd_sc_hd__mux2_1 _10759_ (.A0(\_170_[25] ),
    .A1(\_173_[25] ),
    .S(_04936_),
    .X(_04972_));
 sky130_fd_sc_hd__or2_1 _10760_ (.A(_04971_),
    .B(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__o211a_1 _10761_ (.A1(\_167_[25] ),
    .A2(_04925_),
    .B1(_04973_),
    .C1(_04939_),
    .X(_00594_));
 sky130_fd_sc_hd__or2_1 _10762_ (.A(\_173_[26] ),
    .B(_04953_),
    .X(_04974_));
 sky130_fd_sc_hd__o211a_1 _10763_ (.A1(\_170_[26] ),
    .A2(_04942_),
    .B1(_04958_),
    .C1(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__a211o_1 _10764_ (.A1(\_167_[26] ),
    .A2(_04945_),
    .B1(_04975_),
    .C1(_04952_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _10765_ (.A0(\_170_[27] ),
    .A1(\_173_[27] ),
    .S(_04936_),
    .X(_04976_));
 sky130_fd_sc_hd__or2_1 _10766_ (.A(_04971_),
    .B(_04976_),
    .X(_04977_));
 sky130_fd_sc_hd__o211a_1 _10767_ (.A1(\_167_[27] ),
    .A2(_04925_),
    .B1(_04977_),
    .C1(_04939_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(\_170_[28] ),
    .A1(\_173_[28] ),
    .S(_04936_),
    .X(_04978_));
 sky130_fd_sc_hd__or2_1 _10769_ (.A(_04971_),
    .B(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__o211a_1 _10770_ (.A1(\_167_[28] ),
    .A2(_04925_),
    .B1(_04979_),
    .C1(_04939_),
    .X(_00597_));
 sky130_fd_sc_hd__clkbuf_4 _10771_ (.A(_01225_),
    .X(_04980_));
 sky130_fd_sc_hd__or2_1 _10772_ (.A(\_173_[29] ),
    .B(_04953_),
    .X(_04981_));
 sky130_fd_sc_hd__o211a_1 _10773_ (.A1(\_170_[29] ),
    .A2(_04980_),
    .B1(_04958_),
    .C1(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__a211o_1 _10774_ (.A1(\_167_[29] ),
    .A2(_04945_),
    .B1(_04982_),
    .C1(_04952_),
    .X(_00598_));
 sky130_fd_sc_hd__clkbuf_4 _10775_ (.A(_04671_),
    .X(_04983_));
 sky130_fd_sc_hd__mux2_1 _10776_ (.A0(\_170_[30] ),
    .A1(\_173_[30] ),
    .S(_04936_),
    .X(_04984_));
 sky130_fd_sc_hd__or2_1 _10777_ (.A(_04971_),
    .B(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__o211a_1 _10778_ (.A1(\_167_[30] ),
    .A2(_04983_),
    .B1(_04985_),
    .C1(_04939_),
    .X(_00599_));
 sky130_fd_sc_hd__clkbuf_4 _10779_ (.A(_04682_),
    .X(_04986_));
 sky130_fd_sc_hd__or2_1 _10780_ (.A(\_173_[31] ),
    .B(_04953_),
    .X(_04987_));
 sky130_fd_sc_hd__o211a_1 _10781_ (.A1(\_170_[31] ),
    .A2(_04980_),
    .B1(_04958_),
    .C1(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__a211o_1 _10782_ (.A1(\_167_[31] ),
    .A2(_04986_),
    .B1(_04988_),
    .C1(_04952_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(\_167_[0] ),
    .A1(\_170_[0] ),
    .S(_04936_),
    .X(_04989_));
 sky130_fd_sc_hd__or2_1 _10784_ (.A(_04971_),
    .B(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__o211a_1 _10785_ (.A1(\_164_[0] ),
    .A2(_04983_),
    .B1(_04990_),
    .C1(_04939_),
    .X(_00601_));
 sky130_fd_sc_hd__or2_1 _10786_ (.A(\_170_[1] ),
    .B(_04953_),
    .X(_04991_));
 sky130_fd_sc_hd__o211a_1 _10787_ (.A1(\_167_[1] ),
    .A2(_04980_),
    .B1(_04958_),
    .C1(_04991_),
    .X(_04992_));
 sky130_fd_sc_hd__a211o_1 _10788_ (.A1(\_164_[1] ),
    .A2(_04986_),
    .B1(_04992_),
    .C1(_04952_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(\_167_[2] ),
    .A1(\_170_[2] ),
    .S(_04936_),
    .X(_04993_));
 sky130_fd_sc_hd__or2_1 _10790_ (.A(_04971_),
    .B(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__o211a_1 _10791_ (.A1(\_164_[2] ),
    .A2(_04983_),
    .B1(_04994_),
    .C1(_04939_),
    .X(_00603_));
 sky130_fd_sc_hd__buf_4 _10792_ (.A(_01213_),
    .X(_04995_));
 sky130_fd_sc_hd__mux2_1 _10793_ (.A0(\_167_[3] ),
    .A1(\_170_[3] ),
    .S(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__or2_1 _10794_ (.A(_04971_),
    .B(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__clkbuf_4 _10795_ (.A(_01424_),
    .X(_04998_));
 sky130_fd_sc_hd__o211a_1 _10796_ (.A1(\_164_[3] ),
    .A2(_04983_),
    .B1(_04997_),
    .C1(_04998_),
    .X(_00604_));
 sky130_fd_sc_hd__or2_1 _10797_ (.A(\_170_[4] ),
    .B(_04953_),
    .X(_04999_));
 sky130_fd_sc_hd__o211a_1 _10798_ (.A1(\_167_[4] ),
    .A2(_04980_),
    .B1(_04958_),
    .C1(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__clkbuf_4 _10799_ (.A(_01418_),
    .X(_05001_));
 sky130_fd_sc_hd__a211o_1 _10800_ (.A1(\_164_[4] ),
    .A2(_04986_),
    .B1(_05000_),
    .C1(_05001_),
    .X(_00605_));
 sky130_fd_sc_hd__clkbuf_2 _10801_ (.A(_01216_),
    .X(_05002_));
 sky130_fd_sc_hd__or2_1 _10802_ (.A(\_170_[5] ),
    .B(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__o211a_1 _10803_ (.A1(\_167_[5] ),
    .A2(_04980_),
    .B1(_04958_),
    .C1(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__a211o_1 _10804_ (.A1(\_164_[5] ),
    .A2(_04986_),
    .B1(_05004_),
    .C1(_05001_),
    .X(_00606_));
 sky130_fd_sc_hd__or2_1 _10805_ (.A(\_170_[6] ),
    .B(_05002_),
    .X(_05005_));
 sky130_fd_sc_hd__o211a_1 _10806_ (.A1(\_167_[6] ),
    .A2(_04980_),
    .B1(_04958_),
    .C1(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__a211o_1 _10807_ (.A1(\_164_[6] ),
    .A2(_04986_),
    .B1(_05006_),
    .C1(_05001_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(\_167_[7] ),
    .A1(\_170_[7] ),
    .S(_04995_),
    .X(_05007_));
 sky130_fd_sc_hd__or2_1 _10809_ (.A(_04971_),
    .B(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__o211a_1 _10810_ (.A1(\_164_[7] ),
    .A2(_04983_),
    .B1(_05008_),
    .C1(_04998_),
    .X(_00608_));
 sky130_fd_sc_hd__clkbuf_4 _10811_ (.A(_04685_),
    .X(_05009_));
 sky130_fd_sc_hd__or2_1 _10812_ (.A(\_170_[8] ),
    .B(_05002_),
    .X(_05010_));
 sky130_fd_sc_hd__o211a_1 _10813_ (.A1(\_167_[8] ),
    .A2(_04980_),
    .B1(_05009_),
    .C1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__a211o_1 _10814_ (.A1(\_164_[8] ),
    .A2(_04986_),
    .B1(_05011_),
    .C1(_05001_),
    .X(_00609_));
 sky130_fd_sc_hd__or2_1 _10815_ (.A(\_170_[9] ),
    .B(_05002_),
    .X(_05012_));
 sky130_fd_sc_hd__o211a_1 _10816_ (.A1(\_167_[9] ),
    .A2(_04980_),
    .B1(_05009_),
    .C1(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__a211o_1 _10817_ (.A1(\_164_[9] ),
    .A2(_04986_),
    .B1(_05013_),
    .C1(_05001_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(\_167_[10] ),
    .A1(\_170_[10] ),
    .S(_04995_),
    .X(_05014_));
 sky130_fd_sc_hd__or2_1 _10819_ (.A(_04971_),
    .B(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__o211a_1 _10820_ (.A1(\_164_[10] ),
    .A2(_04983_),
    .B1(_05015_),
    .C1(_04998_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(\_167_[11] ),
    .A1(\_170_[11] ),
    .S(_04995_),
    .X(_05016_));
 sky130_fd_sc_hd__or2_1 _10822_ (.A(_04971_),
    .B(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__o211a_1 _10823_ (.A1(\_164_[11] ),
    .A2(_04983_),
    .B1(_05017_),
    .C1(_04998_),
    .X(_00612_));
 sky130_fd_sc_hd__or2_1 _10824_ (.A(\_170_[12] ),
    .B(_05002_),
    .X(_05018_));
 sky130_fd_sc_hd__o211a_1 _10825_ (.A1(\_167_[12] ),
    .A2(_04980_),
    .B1(_05009_),
    .C1(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__a211o_1 _10826_ (.A1(\_164_[12] ),
    .A2(_04986_),
    .B1(_05019_),
    .C1(_05001_),
    .X(_00613_));
 sky130_fd_sc_hd__or2_1 _10827_ (.A(\_170_[13] ),
    .B(_05002_),
    .X(_05020_));
 sky130_fd_sc_hd__o211a_1 _10828_ (.A1(\_167_[13] ),
    .A2(_04980_),
    .B1(_05009_),
    .C1(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__a211o_1 _10829_ (.A1(\_164_[13] ),
    .A2(_04986_),
    .B1(_05021_),
    .C1(_05001_),
    .X(_00614_));
 sky130_fd_sc_hd__clkbuf_4 _10830_ (.A(_01225_),
    .X(_05022_));
 sky130_fd_sc_hd__or2_1 _10831_ (.A(\_170_[14] ),
    .B(_05002_),
    .X(_05023_));
 sky130_fd_sc_hd__o211a_1 _10832_ (.A1(\_167_[14] ),
    .A2(_05022_),
    .B1(_05009_),
    .C1(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__a211o_1 _10833_ (.A1(\_164_[14] ),
    .A2(_04986_),
    .B1(_05024_),
    .C1(_05001_),
    .X(_00615_));
 sky130_fd_sc_hd__buf_2 _10834_ (.A(_04682_),
    .X(_05025_));
 sky130_fd_sc_hd__or2_1 _10835_ (.A(\_170_[15] ),
    .B(_05002_),
    .X(_05026_));
 sky130_fd_sc_hd__o211a_1 _10836_ (.A1(\_167_[15] ),
    .A2(_05022_),
    .B1(_05009_),
    .C1(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__a211o_1 _10837_ (.A1(\_164_[15] ),
    .A2(_05025_),
    .B1(_05027_),
    .C1(_05001_),
    .X(_00616_));
 sky130_fd_sc_hd__clkbuf_4 _10838_ (.A(_04636_),
    .X(_05028_));
 sky130_fd_sc_hd__mux2_1 _10839_ (.A0(\_167_[16] ),
    .A1(\_170_[16] ),
    .S(_04995_),
    .X(_05029_));
 sky130_fd_sc_hd__or2_1 _10840_ (.A(_05028_),
    .B(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__o211a_1 _10841_ (.A1(\_164_[16] ),
    .A2(_04983_),
    .B1(_05030_),
    .C1(_04998_),
    .X(_00617_));
 sky130_fd_sc_hd__or2_1 _10842_ (.A(\_170_[17] ),
    .B(_05002_),
    .X(_05031_));
 sky130_fd_sc_hd__o211a_1 _10843_ (.A1(\_167_[17] ),
    .A2(_05022_),
    .B1(_05009_),
    .C1(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__a211o_1 _10844_ (.A1(\_164_[17] ),
    .A2(_05025_),
    .B1(_05032_),
    .C1(_05001_),
    .X(_00618_));
 sky130_fd_sc_hd__or2_1 _10845_ (.A(\_170_[18] ),
    .B(_05002_),
    .X(_05033_));
 sky130_fd_sc_hd__o211a_1 _10846_ (.A1(\_167_[18] ),
    .A2(_05022_),
    .B1(_05009_),
    .C1(_05033_),
    .X(_05034_));
 sky130_fd_sc_hd__clkbuf_4 _10847_ (.A(_01418_),
    .X(_05035_));
 sky130_fd_sc_hd__a211o_1 _10848_ (.A1(\_164_[18] ),
    .A2(_05025_),
    .B1(_05034_),
    .C1(_05035_),
    .X(_00619_));
 sky130_fd_sc_hd__clkbuf_2 _10849_ (.A(_01216_),
    .X(_05036_));
 sky130_fd_sc_hd__or2_1 _10850_ (.A(\_170_[19] ),
    .B(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__o211a_1 _10851_ (.A1(\_167_[19] ),
    .A2(_05022_),
    .B1(_05009_),
    .C1(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__a211o_1 _10852_ (.A1(\_164_[19] ),
    .A2(_05025_),
    .B1(_05038_),
    .C1(_05035_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(\_167_[20] ),
    .A1(\_170_[20] ),
    .S(_04995_),
    .X(_05039_));
 sky130_fd_sc_hd__or2_1 _10854_ (.A(_05028_),
    .B(_05039_),
    .X(_05040_));
 sky130_fd_sc_hd__o211a_1 _10855_ (.A1(\_164_[20] ),
    .A2(_04983_),
    .B1(_05040_),
    .C1(_04998_),
    .X(_00621_));
 sky130_fd_sc_hd__or2_1 _10856_ (.A(\_170_[21] ),
    .B(_05036_),
    .X(_05041_));
 sky130_fd_sc_hd__o211a_1 _10857_ (.A1(\_167_[21] ),
    .A2(_05022_),
    .B1(_05009_),
    .C1(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__a211o_1 _10858_ (.A1(\_164_[21] ),
    .A2(_05025_),
    .B1(_05042_),
    .C1(_05035_),
    .X(_00622_));
 sky130_fd_sc_hd__buf_2 _10859_ (.A(_04685_),
    .X(_05043_));
 sky130_fd_sc_hd__or2_1 _10860_ (.A(\_170_[22] ),
    .B(_05036_),
    .X(_05044_));
 sky130_fd_sc_hd__o211a_1 _10861_ (.A1(\_167_[22] ),
    .A2(_05022_),
    .B1(_05043_),
    .C1(_05044_),
    .X(_05045_));
 sky130_fd_sc_hd__a211o_1 _10862_ (.A1(\_164_[22] ),
    .A2(_05025_),
    .B1(_05045_),
    .C1(_05035_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _10863_ (.A0(\_167_[23] ),
    .A1(\_170_[23] ),
    .S(_04995_),
    .X(_05046_));
 sky130_fd_sc_hd__or2_1 _10864_ (.A(_05028_),
    .B(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__o211a_1 _10865_ (.A1(\_164_[23] ),
    .A2(_04983_),
    .B1(_05047_),
    .C1(_04998_),
    .X(_00624_));
 sky130_fd_sc_hd__buf_4 _10866_ (.A(_04671_),
    .X(_05048_));
 sky130_fd_sc_hd__mux2_1 _10867_ (.A0(\_167_[24] ),
    .A1(\_170_[24] ),
    .S(_04995_),
    .X(_05049_));
 sky130_fd_sc_hd__or2_1 _10868_ (.A(_05028_),
    .B(_05049_),
    .X(_05050_));
 sky130_fd_sc_hd__o211a_1 _10869_ (.A1(\_164_[24] ),
    .A2(_05048_),
    .B1(_05050_),
    .C1(_04998_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _10870_ (.A0(\_167_[25] ),
    .A1(\_170_[25] ),
    .S(_04995_),
    .X(_05051_));
 sky130_fd_sc_hd__or2_1 _10871_ (.A(_05028_),
    .B(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__o211a_1 _10872_ (.A1(\_164_[25] ),
    .A2(_05048_),
    .B1(_05052_),
    .C1(_04998_),
    .X(_00626_));
 sky130_fd_sc_hd__or2_1 _10873_ (.A(\_170_[26] ),
    .B(_05036_),
    .X(_05053_));
 sky130_fd_sc_hd__o211a_1 _10874_ (.A1(\_167_[26] ),
    .A2(_05022_),
    .B1(_05043_),
    .C1(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__a211o_1 _10875_ (.A1(\_164_[26] ),
    .A2(_05025_),
    .B1(_05054_),
    .C1(_05035_),
    .X(_00627_));
 sky130_fd_sc_hd__or2_1 _10876_ (.A(\_170_[27] ),
    .B(_05036_),
    .X(_05055_));
 sky130_fd_sc_hd__o211a_1 _10877_ (.A1(\_167_[27] ),
    .A2(_05022_),
    .B1(_05043_),
    .C1(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__a211o_1 _10878_ (.A1(\_164_[27] ),
    .A2(_05025_),
    .B1(_05056_),
    .C1(_05035_),
    .X(_00628_));
 sky130_fd_sc_hd__or2_1 _10879_ (.A(\_170_[28] ),
    .B(_05036_),
    .X(_05057_));
 sky130_fd_sc_hd__o211a_1 _10880_ (.A1(\_167_[28] ),
    .A2(_05022_),
    .B1(_05043_),
    .C1(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__a211o_1 _10881_ (.A1(\_164_[28] ),
    .A2(_05025_),
    .B1(_05058_),
    .C1(_05035_),
    .X(_00629_));
 sky130_fd_sc_hd__clkbuf_4 _10882_ (.A(_01225_),
    .X(_05059_));
 sky130_fd_sc_hd__or2_1 _10883_ (.A(\_170_[29] ),
    .B(_05036_),
    .X(_05060_));
 sky130_fd_sc_hd__o211a_1 _10884_ (.A1(\_167_[29] ),
    .A2(_05059_),
    .B1(_05043_),
    .C1(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__a211o_1 _10885_ (.A1(\_164_[29] ),
    .A2(_05025_),
    .B1(_05061_),
    .C1(_05035_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _10886_ (.A0(\_167_[30] ),
    .A1(\_170_[30] ),
    .S(_04995_),
    .X(_05062_));
 sky130_fd_sc_hd__or2_1 _10887_ (.A(_05028_),
    .B(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__o211a_1 _10888_ (.A1(\_164_[30] ),
    .A2(_05048_),
    .B1(_05063_),
    .C1(_04998_),
    .X(_00631_));
 sky130_fd_sc_hd__buf_4 _10889_ (.A(_01213_),
    .X(_05064_));
 sky130_fd_sc_hd__mux2_1 _10890_ (.A0(\_167_[31] ),
    .A1(\_170_[31] ),
    .S(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__or2_1 _10891_ (.A(_05028_),
    .B(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__clkbuf_4 _10892_ (.A(_01424_),
    .X(_05067_));
 sky130_fd_sc_hd__o211a_1 _10893_ (.A1(\_164_[31] ),
    .A2(_05048_),
    .B1(_05066_),
    .C1(_05067_),
    .X(_00632_));
 sky130_fd_sc_hd__buf_2 _10894_ (.A(_04682_),
    .X(_05068_));
 sky130_fd_sc_hd__or2_1 _10895_ (.A(\_167_[0] ),
    .B(_05036_),
    .X(_05069_));
 sky130_fd_sc_hd__o211a_1 _10896_ (.A1(\_164_[0] ),
    .A2(_05059_),
    .B1(_05043_),
    .C1(_05069_),
    .X(_05070_));
 sky130_fd_sc_hd__a211o_1 _10897_ (.A1(net36),
    .A2(_05068_),
    .B1(_05070_),
    .C1(_05035_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _10898_ (.A0(\_164_[1] ),
    .A1(\_167_[1] ),
    .S(_05064_),
    .X(_05071_));
 sky130_fd_sc_hd__or2_1 _10899_ (.A(_05028_),
    .B(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__o211a_1 _10900_ (.A1(net47),
    .A2(_05048_),
    .B1(_05072_),
    .C1(_05067_),
    .X(_00634_));
 sky130_fd_sc_hd__or2_1 _10901_ (.A(\_167_[2] ),
    .B(_05036_),
    .X(_05073_));
 sky130_fd_sc_hd__o211a_1 _10902_ (.A1(\_164_[2] ),
    .A2(_05059_),
    .B1(_05043_),
    .C1(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__a211o_1 _10903_ (.A1(net58),
    .A2(_05068_),
    .B1(_05074_),
    .C1(_05035_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _10904_ (.A0(\_164_[3] ),
    .A1(\_167_[3] ),
    .S(_05064_),
    .X(_05075_));
 sky130_fd_sc_hd__or2_1 _10905_ (.A(_05028_),
    .B(_05075_),
    .X(_05076_));
 sky130_fd_sc_hd__o211a_1 _10906_ (.A1(net61),
    .A2(_05048_),
    .B1(_05076_),
    .C1(_05067_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(\_164_[4] ),
    .A1(\_167_[4] ),
    .S(_05064_),
    .X(_05077_));
 sky130_fd_sc_hd__or2_1 _10908_ (.A(_05028_),
    .B(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__o211a_1 _10909_ (.A1(net62),
    .A2(_05048_),
    .B1(_05078_),
    .C1(_05067_),
    .X(_00637_));
 sky130_fd_sc_hd__buf_2 _10910_ (.A(_04636_),
    .X(_05079_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(\_164_[5] ),
    .A1(\_167_[5] ),
    .S(_05064_),
    .X(_05080_));
 sky130_fd_sc_hd__or2_1 _10912_ (.A(_05079_),
    .B(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__o211a_1 _10913_ (.A1(net63),
    .A2(_05048_),
    .B1(_05081_),
    .C1(_05067_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _10914_ (.A0(\_164_[6] ),
    .A1(\_167_[6] ),
    .S(_05064_),
    .X(_05082_));
 sky130_fd_sc_hd__or2_1 _10915_ (.A(_05079_),
    .B(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__o211a_1 _10916_ (.A1(net64),
    .A2(_05048_),
    .B1(_05083_),
    .C1(_05067_),
    .X(_00639_));
 sky130_fd_sc_hd__or2_1 _10917_ (.A(\_167_[7] ),
    .B(_05036_),
    .X(_05084_));
 sky130_fd_sc_hd__o211a_1 _10918_ (.A1(\_164_[7] ),
    .A2(_05059_),
    .B1(_05043_),
    .C1(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__buf_2 _10919_ (.A(_01418_),
    .X(_05086_));
 sky130_fd_sc_hd__a211o_1 _10920_ (.A1(net65),
    .A2(_05068_),
    .B1(_05085_),
    .C1(_05086_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _10921_ (.A0(\_164_[8] ),
    .A1(\_167_[8] ),
    .S(_05064_),
    .X(_05087_));
 sky130_fd_sc_hd__or2_1 _10922_ (.A(_05079_),
    .B(_05087_),
    .X(_05088_));
 sky130_fd_sc_hd__o211a_1 _10923_ (.A1(net66),
    .A2(_05048_),
    .B1(_05088_),
    .C1(_05067_),
    .X(_00641_));
 sky130_fd_sc_hd__clkbuf_2 _10924_ (.A(_01216_),
    .X(_05089_));
 sky130_fd_sc_hd__or2_1 _10925_ (.A(\_167_[9] ),
    .B(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__o211a_1 _10926_ (.A1(\_164_[9] ),
    .A2(_05059_),
    .B1(_05043_),
    .C1(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__a211o_1 _10927_ (.A1(net67),
    .A2(_05068_),
    .B1(_05091_),
    .C1(_05086_),
    .X(_00642_));
 sky130_fd_sc_hd__or2_1 _10928_ (.A(\_167_[10] ),
    .B(_05089_),
    .X(_05092_));
 sky130_fd_sc_hd__o211a_1 _10929_ (.A1(\_164_[10] ),
    .A2(_05059_),
    .B1(_05043_),
    .C1(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__a211o_1 _10930_ (.A1(net37),
    .A2(_05068_),
    .B1(_05093_),
    .C1(_05086_),
    .X(_00643_));
 sky130_fd_sc_hd__clkbuf_4 _10931_ (.A(_04685_),
    .X(_05094_));
 sky130_fd_sc_hd__or2_1 _10932_ (.A(\_167_[11] ),
    .B(_05089_),
    .X(_05095_));
 sky130_fd_sc_hd__o211a_1 _10933_ (.A1(\_164_[11] ),
    .A2(_05059_),
    .B1(_05094_),
    .C1(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__a211o_1 _10934_ (.A1(net38),
    .A2(_05068_),
    .B1(_05096_),
    .C1(_05086_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _10935_ (.A0(\_164_[12] ),
    .A1(\_167_[12] ),
    .S(_05064_),
    .X(_05097_));
 sky130_fd_sc_hd__or2_1 _10936_ (.A(_05079_),
    .B(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__o211a_1 _10937_ (.A1(net39),
    .A2(_04853_),
    .B1(_05098_),
    .C1(_05067_),
    .X(_00645_));
 sky130_fd_sc_hd__or2_1 _10938_ (.A(\_167_[13] ),
    .B(_05089_),
    .X(_05099_));
 sky130_fd_sc_hd__o211a_1 _10939_ (.A1(\_164_[13] ),
    .A2(_05059_),
    .B1(_05094_),
    .C1(_05099_),
    .X(_05100_));
 sky130_fd_sc_hd__a211o_1 _10940_ (.A1(net40),
    .A2(_05068_),
    .B1(_05100_),
    .C1(_05086_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _10941_ (.A0(\_164_[14] ),
    .A1(\_167_[14] ),
    .S(_05064_),
    .X(_05101_));
 sky130_fd_sc_hd__or2_1 _10942_ (.A(_05079_),
    .B(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__o211a_1 _10943_ (.A1(net41),
    .A2(_04853_),
    .B1(_05102_),
    .C1(_05067_),
    .X(_00647_));
 sky130_fd_sc_hd__or2_1 _10944_ (.A(\_167_[15] ),
    .B(_05089_),
    .X(_05103_));
 sky130_fd_sc_hd__o211a_1 _10945_ (.A1(\_164_[15] ),
    .A2(_05059_),
    .B1(_05094_),
    .C1(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__a211o_1 _10946_ (.A1(net42),
    .A2(_05068_),
    .B1(_05104_),
    .C1(_05086_),
    .X(_00648_));
 sky130_fd_sc_hd__or2_1 _10947_ (.A(\_167_[16] ),
    .B(_05089_),
    .X(_05105_));
 sky130_fd_sc_hd__o211a_1 _10948_ (.A1(\_164_[16] ),
    .A2(_05059_),
    .B1(_05094_),
    .C1(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__a211o_1 _10949_ (.A1(net43),
    .A2(_05068_),
    .B1(_05106_),
    .C1(_05086_),
    .X(_00649_));
 sky130_fd_sc_hd__clkbuf_4 _10950_ (.A(_01225_),
    .X(_05107_));
 sky130_fd_sc_hd__or2_1 _10951_ (.A(\_167_[17] ),
    .B(_05089_),
    .X(_05108_));
 sky130_fd_sc_hd__o211a_1 _10952_ (.A1(\_164_[17] ),
    .A2(_05107_),
    .B1(_05094_),
    .C1(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__a211o_1 _10953_ (.A1(net44),
    .A2(_05068_),
    .B1(_05109_),
    .C1(_05086_),
    .X(_00650_));
 sky130_fd_sc_hd__clkbuf_4 _10954_ (.A(_04682_),
    .X(_05110_));
 sky130_fd_sc_hd__or2_1 _10955_ (.A(\_167_[18] ),
    .B(_05089_),
    .X(_05111_));
 sky130_fd_sc_hd__o211a_1 _10956_ (.A1(\_164_[18] ),
    .A2(_05107_),
    .B1(_05094_),
    .C1(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__a211o_1 _10957_ (.A1(net45),
    .A2(_05110_),
    .B1(_05112_),
    .C1(_05086_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _10958_ (.A0(\_164_[19] ),
    .A1(\_167_[19] ),
    .S(_05064_),
    .X(_05113_));
 sky130_fd_sc_hd__or2_1 _10959_ (.A(_05079_),
    .B(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__o211a_1 _10960_ (.A1(net46),
    .A2(_04853_),
    .B1(_05114_),
    .C1(_05067_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _10961_ (.A0(\_164_[20] ),
    .A1(\_167_[20] ),
    .S(_01214_),
    .X(_05115_));
 sky130_fd_sc_hd__or2_1 _10962_ (.A(_05079_),
    .B(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__buf_2 _10963_ (.A(_01424_),
    .X(_05117_));
 sky130_fd_sc_hd__o211a_1 _10964_ (.A1(net48),
    .A2(_04853_),
    .B1(_05116_),
    .C1(_05117_),
    .X(_00653_));
 sky130_fd_sc_hd__or2_1 _10965_ (.A(\_167_[21] ),
    .B(_05089_),
    .X(_05118_));
 sky130_fd_sc_hd__o211a_1 _10966_ (.A1(\_164_[21] ),
    .A2(_05107_),
    .B1(_05094_),
    .C1(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__a211o_1 _10967_ (.A1(net49),
    .A2(_05110_),
    .B1(_05119_),
    .C1(_05086_),
    .X(_00654_));
 sky130_fd_sc_hd__or2_1 _10968_ (.A(\_167_[22] ),
    .B(_05089_),
    .X(_05120_));
 sky130_fd_sc_hd__o211a_1 _10969_ (.A1(\_164_[22] ),
    .A2(_05107_),
    .B1(_05094_),
    .C1(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__buf_4 _10970_ (.A(_01435_),
    .X(_05122_));
 sky130_fd_sc_hd__a211o_1 _10971_ (.A1(net50),
    .A2(_05110_),
    .B1(_05121_),
    .C1(_05122_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _10972_ (.A0(\_164_[23] ),
    .A1(\_167_[23] ),
    .S(_01214_),
    .X(_05123_));
 sky130_fd_sc_hd__or2_1 _10973_ (.A(_05079_),
    .B(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__o211a_1 _10974_ (.A1(net51),
    .A2(_04853_),
    .B1(_05124_),
    .C1(_05117_),
    .X(_00656_));
 sky130_fd_sc_hd__or2_1 _10975_ (.A(\_167_[24] ),
    .B(_04867_),
    .X(_05125_));
 sky130_fd_sc_hd__o211a_1 _10976_ (.A1(\_164_[24] ),
    .A2(_05107_),
    .B1(_05094_),
    .C1(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__a211o_1 _10977_ (.A1(net52),
    .A2(_05110_),
    .B1(_05126_),
    .C1(_05122_),
    .X(_00657_));
 sky130_fd_sc_hd__or2_1 _10978_ (.A(\_167_[25] ),
    .B(_04867_),
    .X(_05127_));
 sky130_fd_sc_hd__o211a_1 _10979_ (.A1(\_164_[25] ),
    .A2(_05107_),
    .B1(_05094_),
    .C1(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__a211o_1 _10980_ (.A1(net53),
    .A2(_05110_),
    .B1(_05128_),
    .C1(_05122_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _10981_ (.A0(\_164_[26] ),
    .A1(\_167_[26] ),
    .S(_01214_),
    .X(_05129_));
 sky130_fd_sc_hd__or2_1 _10982_ (.A(_05079_),
    .B(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__o211a_1 _10983_ (.A1(net54),
    .A2(_04853_),
    .B1(_05130_),
    .C1(_05117_),
    .X(_00659_));
 sky130_fd_sc_hd__or2_1 _10984_ (.A(\_167_[27] ),
    .B(_04867_),
    .X(_05131_));
 sky130_fd_sc_hd__o211a_1 _10985_ (.A1(\_164_[27] ),
    .A2(_05107_),
    .B1(_04865_),
    .C1(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__a211o_1 _10986_ (.A1(net55),
    .A2(_05110_),
    .B1(_05132_),
    .C1(_05122_),
    .X(_00660_));
 sky130_fd_sc_hd__or2_1 _10987_ (.A(\_167_[28] ),
    .B(_04867_),
    .X(_05133_));
 sky130_fd_sc_hd__o211a_1 _10988_ (.A1(\_164_[28] ),
    .A2(_05107_),
    .B1(_04865_),
    .C1(_05133_),
    .X(_05134_));
 sky130_fd_sc_hd__a211o_1 _10989_ (.A1(net56),
    .A2(_05110_),
    .B1(_05134_),
    .C1(_05122_),
    .X(_00661_));
 sky130_fd_sc_hd__or2_1 _10990_ (.A(\_167_[29] ),
    .B(_04867_),
    .X(_05135_));
 sky130_fd_sc_hd__o211a_1 _10991_ (.A1(\_164_[29] ),
    .A2(_05107_),
    .B1(_04865_),
    .C1(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__a211o_1 _10992_ (.A1(net57),
    .A2(_05110_),
    .B1(_05136_),
    .C1(_05122_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _10993_ (.A0(\_164_[30] ),
    .A1(\_167_[30] ),
    .S(_01214_),
    .X(_05137_));
 sky130_fd_sc_hd__or2_1 _10994_ (.A(_05079_),
    .B(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__o211a_1 _10995_ (.A1(net59),
    .A2(_04853_),
    .B1(_05138_),
    .C1(_05117_),
    .X(_00663_));
 sky130_fd_sc_hd__or2_1 _10996_ (.A(\_167_[31] ),
    .B(_04867_),
    .X(_05139_));
 sky130_fd_sc_hd__o211a_1 _10997_ (.A1(\_164_[31] ),
    .A2(_05107_),
    .B1(_04865_),
    .C1(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__a211o_1 _10998_ (.A1(net60),
    .A2(_05110_),
    .B1(_05140_),
    .C1(_05122_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _10999_ (.A0(net36),
    .A1(\_164_[0] ),
    .S(_01215_),
    .X(_05141_));
 sky130_fd_sc_hd__nor2_1 _11000_ (.A(_02886_),
    .B(_04631_),
    .Y(_05142_));
 sky130_fd_sc_hd__a211o_1 _11001_ (.A1(_04855_),
    .A2(_05141_),
    .B1(_05142_),
    .C1(_05122_),
    .X(_00665_));
 sky130_fd_sc_hd__a221o_1 _11002_ (.A1(\_164_[1] ),
    .A2(net68),
    .B1(_02907_),
    .B2(_04692_),
    .C1(_02711_),
    .X(_05143_));
 sky130_fd_sc_hd__a21o_1 _11003_ (.A1(net47),
    .A2(_04849_),
    .B1(_05143_),
    .X(_00666_));
 sky130_fd_sc_hd__a221o_1 _11004_ (.A1(\_164_[2] ),
    .A2(net68),
    .B1(_02936_),
    .B2(_04692_),
    .C1(_01417_),
    .X(_05144_));
 sky130_fd_sc_hd__a21o_1 _11005_ (.A1(net58),
    .A2(_04849_),
    .B1(_05144_),
    .X(_00667_));
 sky130_fd_sc_hd__o221a_1 _11006_ (.A1(\_164_[3] ),
    .A2(_04678_),
    .B1(_02946_),
    .B2(_04686_),
    .C1(_04648_),
    .X(_05145_));
 sky130_fd_sc_hd__o21a_1 _11007_ (.A1(net61),
    .A2(_04629_),
    .B1(_05145_),
    .X(_00668_));
 sky130_fd_sc_hd__o221a_1 _11008_ (.A1(\_164_[4] ),
    .A2(_04678_),
    .B1(_02977_),
    .B2(_04686_),
    .C1(_04648_),
    .X(_05146_));
 sky130_fd_sc_hd__o21a_1 _11009_ (.A1(net62),
    .A2(_04629_),
    .B1(_05146_),
    .X(_00669_));
 sky130_fd_sc_hd__a221o_1 _11010_ (.A1(\_164_[5] ),
    .A2(net68),
    .B1(_03030_),
    .B2(_04692_),
    .C1(_01417_),
    .X(_05147_));
 sky130_fd_sc_hd__a21o_1 _11011_ (.A1(net63),
    .A2(_04849_),
    .B1(_05147_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _11012_ (.A0(net64),
    .A1(\_164_[6] ),
    .S(_01215_),
    .X(_05148_));
 sky130_fd_sc_hd__nor2_1 _11013_ (.A(_03060_),
    .B(_04631_),
    .Y(_05149_));
 sky130_fd_sc_hd__a211o_1 _11014_ (.A1(_04855_),
    .A2(_05148_),
    .B1(_05149_),
    .C1(_05122_),
    .X(_00671_));
 sky130_fd_sc_hd__o221a_1 _11015_ (.A1(\_164_[7] ),
    .A2(_04678_),
    .B1(_03069_),
    .B2(_04686_),
    .C1(_04648_),
    .X(_05150_));
 sky130_fd_sc_hd__o21a_1 _11016_ (.A1(net65),
    .A2(_04629_),
    .B1(_05150_),
    .X(_00672_));
 sky130_fd_sc_hd__o2bb2a_1 _11017_ (.A1_N(_03125_),
    .A2_N(_04682_),
    .B1(_04627_),
    .B2(net66),
    .X(_05151_));
 sky130_fd_sc_hd__o211a_1 _11018_ (.A1(\_164_[8] ),
    .A2(_01218_),
    .B1(_03864_),
    .C1(_05151_),
    .X(_00673_));
 sky130_fd_sc_hd__a221o_1 _11019_ (.A1(\_164_[9] ),
    .A2(net68),
    .B1(_03133_),
    .B2(_04692_),
    .C1(_01417_),
    .X(_05152_));
 sky130_fd_sc_hd__a21o_1 _11020_ (.A1(net67),
    .A2(_04849_),
    .B1(_05152_),
    .X(_00674_));
 sky130_fd_sc_hd__a2bb2o_1 _11021_ (.A1_N(_03184_),
    .A2_N(_04865_),
    .B1(\_164_[10] ),
    .B2(_04684_),
    .X(_05153_));
 sky130_fd_sc_hd__a211o_1 _11022_ (.A1(net37),
    .A2(_04848_),
    .B1(_05153_),
    .C1(_05122_),
    .X(_00675_));
 sky130_fd_sc_hd__nor2_1 _11023_ (.A(_03215_),
    .B(_04630_),
    .Y(_05154_));
 sky130_fd_sc_hd__a211o_1 _11024_ (.A1(\_164_[11] ),
    .A2(_04865_),
    .B1(_04638_),
    .C1(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__o211a_1 _11025_ (.A1(net38),
    .A2(_04628_),
    .B1(_05155_),
    .C1(_05117_),
    .X(_00676_));
 sky130_fd_sc_hd__o221a_1 _11026_ (.A1(\_164_[12] ),
    .A2(_01217_),
    .B1(_04627_),
    .B2(net39),
    .C1(_02833_),
    .X(_05156_));
 sky130_fd_sc_hd__a21boi_1 _11027_ (.A1(_03248_),
    .A2(_04861_),
    .B1_N(_05156_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _11028_ (.A(_03275_),
    .B(_04636_),
    .Y(_05157_));
 sky130_fd_sc_hd__o221a_1 _11029_ (.A1(\_164_[13] ),
    .A2(_01217_),
    .B1(_04627_),
    .B2(net40),
    .C1(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__or2_1 _11030_ (.A(_01710_),
    .B(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__clkbuf_1 _11031_ (.A(_05159_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(net41),
    .A1(\_164_[14] ),
    .S(_01215_),
    .X(_05160_));
 sky130_fd_sc_hd__nor2_1 _11033_ (.A(_03306_),
    .B(_04631_),
    .Y(_05161_));
 sky130_fd_sc_hd__a211o_1 _11034_ (.A1(_04855_),
    .A2(_05160_),
    .B1(_05161_),
    .C1(_01436_),
    .X(_00679_));
 sky130_fd_sc_hd__nand2_1 _11035_ (.A(_03338_),
    .B(_04681_),
    .Y(_05162_));
 sky130_fd_sc_hd__o211a_1 _11036_ (.A1(\_164_[15] ),
    .A2(_04872_),
    .B1(_04633_),
    .C1(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__a211o_1 _11037_ (.A1(net42),
    .A2(_04848_),
    .B1(_05163_),
    .C1(_01436_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _11038_ (.A0(net43),
    .A1(\_164_[16] ),
    .S(_01215_),
    .X(_05164_));
 sky130_fd_sc_hd__nor2_1 _11039_ (.A(_03376_),
    .B(_04631_),
    .Y(_05165_));
 sky130_fd_sc_hd__a211o_1 _11040_ (.A1(_04855_),
    .A2(_05164_),
    .B1(_05165_),
    .C1(_01436_),
    .X(_00681_));
 sky130_fd_sc_hd__nor2_1 _11041_ (.A(_03407_),
    .B(_04630_),
    .Y(_05166_));
 sky130_fd_sc_hd__a211o_1 _11042_ (.A1(\_164_[17] ),
    .A2(_04865_),
    .B1(_04638_),
    .C1(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__o211a_1 _11043_ (.A1(net44),
    .A2(_04628_),
    .B1(_05167_),
    .C1(_05117_),
    .X(_00682_));
 sky130_fd_sc_hd__o221a_1 _11044_ (.A1(\_164_[18] ),
    .A2(_01217_),
    .B1(_04627_),
    .B2(net45),
    .C1(_02833_),
    .X(_05168_));
 sky130_fd_sc_hd__a21boi_1 _11045_ (.A1(_03438_),
    .A2(_04861_),
    .B1_N(_05168_),
    .Y(_00683_));
 sky130_fd_sc_hd__nand2_1 _11046_ (.A(_03464_),
    .B(_04681_),
    .Y(_05169_));
 sky130_fd_sc_hd__o211a_1 _11047_ (.A1(\_164_[19] ),
    .A2(_04872_),
    .B1(_04633_),
    .C1(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__a211o_1 _11048_ (.A1(net46),
    .A2(_04848_),
    .B1(_05170_),
    .C1(_01436_),
    .X(_00684_));
 sky130_fd_sc_hd__o21a_1 _11049_ (.A1(\_164_[20] ),
    .A2(_01218_),
    .B1(_04648_),
    .X(_05171_));
 sky130_fd_sc_hd__o221a_1 _11050_ (.A1(_03478_),
    .A2(_04855_),
    .B1(_04628_),
    .B2(net48),
    .C1(_05171_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _11051_ (.A0(\_164_[21] ),
    .A1(_03512_),
    .S(_04636_),
    .X(_05172_));
 sky130_fd_sc_hd__or2_1 _11052_ (.A(_04638_),
    .B(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__o211a_1 _11053_ (.A1(net49),
    .A2(_04628_),
    .B1(_05173_),
    .C1(_05117_),
    .X(_00686_));
 sky130_fd_sc_hd__o221a_1 _11054_ (.A1(\_164_[22] ),
    .A2(_01217_),
    .B1(_04627_),
    .B2(net50),
    .C1(_01423_),
    .X(_05174_));
 sky130_fd_sc_hd__a21boi_1 _11055_ (.A1(_03544_),
    .A2(_04861_),
    .B1_N(_05174_),
    .Y(_00687_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(\_164_[23] ),
    .A1(_03595_),
    .S(_04636_),
    .X(_05175_));
 sky130_fd_sc_hd__or2_1 _11057_ (.A(_04638_),
    .B(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__o211a_1 _11058_ (.A1(net51),
    .A2(_04628_),
    .B1(_05176_),
    .C1(_05117_),
    .X(_00688_));
 sky130_fd_sc_hd__o21a_1 _11059_ (.A1(\_164_[24] ),
    .A2(_01218_),
    .B1(_04648_),
    .X(_05177_));
 sky130_fd_sc_hd__o221a_1 _11060_ (.A1(_03607_),
    .A2(_04855_),
    .B1(_04628_),
    .B2(net52),
    .C1(_05177_),
    .X(_00689_));
 sky130_fd_sc_hd__or2_1 _11061_ (.A(\_164_[25] ),
    .B(_04867_),
    .X(_05178_));
 sky130_fd_sc_hd__o211a_1 _11062_ (.A1(net53),
    .A2(_01226_),
    .B1(_04865_),
    .C1(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__a211o_1 _11063_ (.A1(_03667_),
    .A2(_05110_),
    .B1(_05179_),
    .C1(_01436_),
    .X(_00690_));
 sky130_fd_sc_hd__o21a_1 _11064_ (.A1(\_164_[26] ),
    .A2(_01218_),
    .B1(_04648_),
    .X(_05180_));
 sky130_fd_sc_hd__o221a_1 _11065_ (.A1(_03704_),
    .A2(_04855_),
    .B1(_04628_),
    .B2(net54),
    .C1(_05180_),
    .X(_00691_));
 sky130_fd_sc_hd__nand2_1 _11066_ (.A(_03735_),
    .B(_04681_),
    .Y(_05181_));
 sky130_fd_sc_hd__o211a_1 _11067_ (.A1(\_164_[27] ),
    .A2(_04872_),
    .B1(_04633_),
    .C1(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__a211o_1 _11068_ (.A1(net55),
    .A2(_04848_),
    .B1(_05182_),
    .C1(_01436_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _11069_ (.A0(\_164_[28] ),
    .A1(_03774_),
    .S(_04636_),
    .X(_05183_));
 sky130_fd_sc_hd__or2_1 _11070_ (.A(_04638_),
    .B(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__o211a_1 _11071_ (.A1(net56),
    .A2(_04628_),
    .B1(_05184_),
    .C1(_05117_),
    .X(_00693_));
 sky130_fd_sc_hd__or2_1 _11072_ (.A(_03810_),
    .B(_04625_),
    .X(_05185_));
 sky130_fd_sc_hd__o211a_1 _11073_ (.A1(\_164_[29] ),
    .A2(_04872_),
    .B1(_04627_),
    .C1(_05185_),
    .X(_05186_));
 sky130_fd_sc_hd__a211o_1 _11074_ (.A1(net57),
    .A2(_04848_),
    .B1(_05186_),
    .C1(_01436_),
    .X(_00694_));
 sky130_fd_sc_hd__a221o_1 _11075_ (.A1(\_164_[30] ),
    .A2(_01226_),
    .B1(_04637_),
    .B2(net59),
    .C1(_01417_),
    .X(_05187_));
 sky130_fd_sc_hd__o21bai_1 _11076_ (.A1(_03841_),
    .A2(_04691_),
    .B1_N(_05187_),
    .Y(_00695_));
 sky130_fd_sc_hd__o21a_1 _11077_ (.A1(\_164_[31] ),
    .A2(_01217_),
    .B1(_04630_),
    .X(_05188_));
 sky130_fd_sc_hd__a21o_1 _11078_ (.A1(_03862_),
    .A2(_04724_),
    .B1(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__o211a_1 _11079_ (.A1(net60),
    .A2(_04628_),
    .B1(_05189_),
    .C1(_05117_),
    .X(_00696_));
 sky130_fd_sc_hd__inv_2 _11080_ (.A(_03866_),
    .Y(_00111_));
 sky130_fd_sc_hd__inv_2 _11081_ (.A(_03866_),
    .Y(_00112_));
 sky130_fd_sc_hd__inv_2 _11082_ (.A(_03866_),
    .Y(_00113_));
 sky130_fd_sc_hd__inv_2 _11083_ (.A(_03866_),
    .Y(_00114_));
 sky130_fd_sc_hd__nor2_4 _11084_ (.A(net35),
    .B(_01325_),
    .Y(_05190_));
 sky130_fd_sc_hd__nor2_4 _11085_ (.A(net35),
    .B(_01248_),
    .Y(_05191_));
 sky130_fd_sc_hd__nor2_4 _11086_ (.A(_05190_),
    .B(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__clkbuf_4 _11087_ (.A(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__nand2_4 _11088_ (.A(_01303_),
    .B(_01318_),
    .Y(_05194_));
 sky130_fd_sc_hd__or2_1 _11089_ (.A(net35),
    .B(_01325_),
    .X(_05195_));
 sky130_fd_sc_hd__buf_2 _11090_ (.A(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__o21ai_1 _11091_ (.A1(\_158_[0] ),
    .A2(_05194_),
    .B1(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__or2_1 _11092_ (.A(net32),
    .B(_05196_),
    .X(_05198_));
 sky130_fd_sc_hd__a22o_1 _11093_ (.A1(\_158_[0] ),
    .A2(_05193_),
    .B1(_05197_),
    .B2(_05198_),
    .X(_00701_));
 sky130_fd_sc_hd__inv_2 _11094_ (.A(\_158_[1] ),
    .Y(_05199_));
 sky130_fd_sc_hd__nor2_1 _11095_ (.A(net2),
    .B(_05196_),
    .Y(_05200_));
 sky130_fd_sc_hd__o31a_1 _11096_ (.A1(\_158_[1] ),
    .A2(\_158_[0] ),
    .A3(_05194_),
    .B1(_05196_),
    .X(_05201_));
 sky130_fd_sc_hd__o22ai_1 _11097_ (.A1(_05199_),
    .A2(_05197_),
    .B1(_05200_),
    .B2(_05201_),
    .Y(_00702_));
 sky130_fd_sc_hd__buf_2 _11098_ (.A(_05190_),
    .X(_05202_));
 sky130_fd_sc_hd__nor3_1 _11099_ (.A(\_158_[1] ),
    .B(\_158_[0] ),
    .C(\_158_[2] ),
    .Y(_05203_));
 sky130_fd_sc_hd__o311a_1 _11100_ (.A1(\_158_[1] ),
    .A2(\_158_[0] ),
    .A3(_05194_),
    .B1(_05196_),
    .C1(\_158_[2] ),
    .X(_05204_));
 sky130_fd_sc_hd__a221o_1 _11101_ (.A1(net3),
    .A2(_05202_),
    .B1(_05191_),
    .B2(_05203_),
    .C1(_05204_),
    .X(_00703_));
 sky130_fd_sc_hd__or2b_1 _11102_ (.A(_05203_),
    .B_N(\_158_[3] ),
    .X(_05205_));
 sky130_fd_sc_hd__a21oi_1 _11103_ (.A1(_01254_),
    .A2(_05205_),
    .B1(_05194_),
    .Y(_05206_));
 sky130_fd_sc_hd__a221o_1 _11104_ (.A1(net4),
    .A2(_05202_),
    .B1(_05193_),
    .B2(\_158_[3] ),
    .C1(_05206_),
    .X(_00704_));
 sky130_fd_sc_hd__nor2_1 _11105_ (.A(net5),
    .B(_05196_),
    .Y(_05207_));
 sky130_fd_sc_hd__o31a_1 _11106_ (.A1(\_158_[4] ),
    .A2(_01254_),
    .A3(_05194_),
    .B1(_05196_),
    .X(_05208_));
 sky130_fd_sc_hd__o211ai_1 _11107_ (.A1(_01254_),
    .A2(_05194_),
    .B1(_05196_),
    .C1(\_158_[4] ),
    .Y(_05209_));
 sky130_fd_sc_hd__o21ai_1 _11108_ (.A1(_05207_),
    .A2(_05208_),
    .B1(_05209_),
    .Y(_00705_));
 sky130_fd_sc_hd__o21ai_1 _11109_ (.A1(\_158_[4] ),
    .A2(_01254_),
    .B1(\_158_[5] ),
    .Y(_05210_));
 sky130_fd_sc_hd__nand2_1 _11110_ (.A(_01255_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__mux2_1 _11111_ (.A0(net6),
    .A1(_05211_),
    .S(_05196_),
    .X(_05212_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(_05212_),
    .A1(\_158_[5] ),
    .S(_05192_),
    .X(_05213_));
 sky130_fd_sc_hd__clkbuf_1 _11113_ (.A(_05213_),
    .X(_00706_));
 sky130_fd_sc_hd__nand2_1 _11114_ (.A(\_158_[6] ),
    .B(_01255_),
    .Y(_05214_));
 sky130_fd_sc_hd__nand2_1 _11115_ (.A(_01256_),
    .B(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__mux2_1 _11116_ (.A0(net7),
    .A1(_05215_),
    .S(_05195_),
    .X(_05216_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(_05216_),
    .A1(\_158_[6] ),
    .S(_05192_),
    .X(_05217_));
 sky130_fd_sc_hd__clkbuf_1 _11118_ (.A(_05217_),
    .X(_00707_));
 sky130_fd_sc_hd__xnor2_1 _11119_ (.A(\_158_[7] ),
    .B(_01256_),
    .Y(_05218_));
 sky130_fd_sc_hd__and2_1 _11120_ (.A(net8),
    .B(_05190_),
    .X(_05219_));
 sky130_fd_sc_hd__a221o_1 _11121_ (.A1(\_158_[7] ),
    .A2(_05193_),
    .B1(_05218_),
    .B2(_05191_),
    .C1(_05219_),
    .X(_00708_));
 sky130_fd_sc_hd__o21ai_1 _11122_ (.A1(\_158_[7] ),
    .A2(_01256_),
    .B1(\_158_[8] ),
    .Y(_05220_));
 sky130_fd_sc_hd__nand2_1 _11123_ (.A(_01257_),
    .B(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__and2_1 _11124_ (.A(net9),
    .B(_05190_),
    .X(_05222_));
 sky130_fd_sc_hd__a221o_1 _11125_ (.A1(\_158_[8] ),
    .A2(_05193_),
    .B1(_05221_),
    .B2(_05191_),
    .C1(_05222_),
    .X(_00709_));
 sky130_fd_sc_hd__nand2_1 _11126_ (.A(\_158_[9] ),
    .B(_01257_),
    .Y(_05223_));
 sky130_fd_sc_hd__a21oi_1 _11127_ (.A1(_01258_),
    .A2(_05223_),
    .B1(_05194_),
    .Y(_05224_));
 sky130_fd_sc_hd__a22o_1 _11128_ (.A1(net10),
    .A2(_05190_),
    .B1(_05192_),
    .B2(\_158_[9] ),
    .X(_05225_));
 sky130_fd_sc_hd__or2_1 _11129_ (.A(_05224_),
    .B(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__clkbuf_1 _11130_ (.A(_05226_),
    .X(_00710_));
 sky130_fd_sc_hd__clkbuf_4 _11131_ (.A(_05191_),
    .X(_05227_));
 sky130_fd_sc_hd__xnor2_1 _11132_ (.A(\_158_[10] ),
    .B(_01258_),
    .Y(_05228_));
 sky130_fd_sc_hd__a22o_1 _11133_ (.A1(net11),
    .A2(_05202_),
    .B1(_05193_),
    .B2(\_158_[10] ),
    .X(_05229_));
 sky130_fd_sc_hd__a21o_1 _11134_ (.A1(_05227_),
    .A2(_05228_),
    .B1(_05229_),
    .X(_00711_));
 sky130_fd_sc_hd__o21ai_1 _11135_ (.A1(\_158_[10] ),
    .A2(_01258_),
    .B1(\_158_[11] ),
    .Y(_05230_));
 sky130_fd_sc_hd__nand2_1 _11136_ (.A(_01259_),
    .B(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__a22o_1 _11137_ (.A1(net13),
    .A2(_05202_),
    .B1(_05193_),
    .B2(\_158_[11] ),
    .X(_05232_));
 sky130_fd_sc_hd__a21o_1 _11138_ (.A1(_05227_),
    .A2(_05231_),
    .B1(_05232_),
    .X(_00712_));
 sky130_fd_sc_hd__nand2_1 _11139_ (.A(\_158_[12] ),
    .B(_01259_),
    .Y(_05233_));
 sky130_fd_sc_hd__a21oi_1 _11140_ (.A1(_01260_),
    .A2(_05233_),
    .B1(_05194_),
    .Y(_05234_));
 sky130_fd_sc_hd__a22o_1 _11141_ (.A1(net14),
    .A2(_05190_),
    .B1(_05192_),
    .B2(\_158_[12] ),
    .X(_05235_));
 sky130_fd_sc_hd__or2_1 _11142_ (.A(_05234_),
    .B(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__clkbuf_1 _11143_ (.A(_05236_),
    .X(_00713_));
 sky130_fd_sc_hd__xnor2_1 _11144_ (.A(\_158_[13] ),
    .B(_01260_),
    .Y(_05237_));
 sky130_fd_sc_hd__a22o_1 _11145_ (.A1(net15),
    .A2(_05202_),
    .B1(_05193_),
    .B2(\_158_[13] ),
    .X(_05238_));
 sky130_fd_sc_hd__a21o_1 _11146_ (.A1(_05227_),
    .A2(_05237_),
    .B1(_05238_),
    .X(_00714_));
 sky130_fd_sc_hd__o21ai_1 _11147_ (.A1(\_158_[13] ),
    .A2(_01260_),
    .B1(\_158_[14] ),
    .Y(_05239_));
 sky130_fd_sc_hd__nand2_1 _11148_ (.A(_01261_),
    .B(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__a22o_1 _11149_ (.A1(net16),
    .A2(_05202_),
    .B1(_05193_),
    .B2(\_158_[14] ),
    .X(_05241_));
 sky130_fd_sc_hd__a21o_1 _11150_ (.A1(_05227_),
    .A2(_05240_),
    .B1(_05241_),
    .X(_00715_));
 sky130_fd_sc_hd__nand2_1 _11151_ (.A(\_158_[15] ),
    .B(_01261_),
    .Y(_05242_));
 sky130_fd_sc_hd__a21oi_1 _11152_ (.A1(_01262_),
    .A2(_05242_),
    .B1(_05194_),
    .Y(_05243_));
 sky130_fd_sc_hd__a22o_1 _11153_ (.A1(net17),
    .A2(_05190_),
    .B1(_05192_),
    .B2(\_158_[15] ),
    .X(_05244_));
 sky130_fd_sc_hd__or2_1 _11154_ (.A(_05243_),
    .B(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__clkbuf_1 _11155_ (.A(_05245_),
    .X(_00716_));
 sky130_fd_sc_hd__xnor2_1 _11156_ (.A(\_158_[16] ),
    .B(_01262_),
    .Y(_05246_));
 sky130_fd_sc_hd__a22o_1 _11157_ (.A1(net18),
    .A2(_05202_),
    .B1(_05193_),
    .B2(\_158_[16] ),
    .X(_05247_));
 sky130_fd_sc_hd__a21o_1 _11158_ (.A1(_05227_),
    .A2(_05246_),
    .B1(_05247_),
    .X(_00717_));
 sky130_fd_sc_hd__o21ai_1 _11159_ (.A1(\_158_[16] ),
    .A2(_01262_),
    .B1(\_158_[17] ),
    .Y(_05248_));
 sky130_fd_sc_hd__nand2_1 _11160_ (.A(_01263_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__a22o_1 _11161_ (.A1(net19),
    .A2(_05202_),
    .B1(_05193_),
    .B2(\_158_[17] ),
    .X(_05250_));
 sky130_fd_sc_hd__a21o_1 _11162_ (.A1(_05227_),
    .A2(_05249_),
    .B1(_05250_),
    .X(_00718_));
 sky130_fd_sc_hd__nand2_1 _11163_ (.A(\_158_[18] ),
    .B(_01263_),
    .Y(_05251_));
 sky130_fd_sc_hd__nand2_1 _11164_ (.A(_01264_),
    .B(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hd__a22o_1 _11165_ (.A1(net20),
    .A2(_05202_),
    .B1(_05192_),
    .B2(\_158_[18] ),
    .X(_05253_));
 sky130_fd_sc_hd__a21o_1 _11166_ (.A1(_05227_),
    .A2(_05252_),
    .B1(_05253_),
    .X(_00719_));
 sky130_fd_sc_hd__xnor2_1 _11167_ (.A(\_158_[19] ),
    .B(_01264_),
    .Y(_05254_));
 sky130_fd_sc_hd__a22o_1 _11168_ (.A1(net21),
    .A2(_05202_),
    .B1(_05192_),
    .B2(\_158_[19] ),
    .X(_05255_));
 sky130_fd_sc_hd__a21o_1 _11169_ (.A1(_05227_),
    .A2(_05254_),
    .B1(_05255_),
    .X(_00720_));
 sky130_fd_sc_hd__o21ai_1 _11170_ (.A1(\_158_[19] ),
    .A2(_01264_),
    .B1(\_158_[20] ),
    .Y(_05256_));
 sky130_fd_sc_hd__nand2_1 _11171_ (.A(_01265_),
    .B(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__a22o_1 _11172_ (.A1(net22),
    .A2(_05190_),
    .B1(_05192_),
    .B2(\_158_[20] ),
    .X(_05258_));
 sky130_fd_sc_hd__a21o_1 _11173_ (.A1(_05227_),
    .A2(_05257_),
    .B1(_05258_),
    .X(_00721_));
 sky130_fd_sc_hd__nand2_1 _11174_ (.A(\_158_[21] ),
    .B(_01265_),
    .Y(_05259_));
 sky130_fd_sc_hd__nand2_1 _11175_ (.A(_01266_),
    .B(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__a22o_1 _11176_ (.A1(net24),
    .A2(_05190_),
    .B1(_05192_),
    .B2(\_158_[21] ),
    .X(_05261_));
 sky130_fd_sc_hd__a21o_1 _11177_ (.A1(_05227_),
    .A2(_05260_),
    .B1(_05261_),
    .X(_00722_));
 sky130_fd_sc_hd__clkbuf_4 _11178_ (.A(_01368_),
    .X(_05262_));
 sky130_fd_sc_hd__clkbuf_4 _11179_ (.A(_01361_),
    .X(_05263_));
 sky130_fd_sc_hd__nand2_1 _11180_ (.A(\_149_[0] ),
    .B(\_132_[0] ),
    .Y(_05264_));
 sky130_fd_sc_hd__or2_1 _11181_ (.A(\_149_[0] ),
    .B(\_132_[0] ),
    .X(_05265_));
 sky130_fd_sc_hd__and3_1 _11182_ (.A(_05263_),
    .B(_05264_),
    .C(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__a21o_1 _11183_ (.A1(\_152_[0] ),
    .A2(_05262_),
    .B1(_05266_),
    .X(_00723_));
 sky130_fd_sc_hd__and2_1 _11184_ (.A(\_149_[1] ),
    .B(\_132_[1] ),
    .X(_05267_));
 sky130_fd_sc_hd__nor2_1 _11185_ (.A(\_149_[1] ),
    .B(\_132_[1] ),
    .Y(_05268_));
 sky130_fd_sc_hd__nor2_1 _11186_ (.A(_05267_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__xnor2_1 _11187_ (.A(_05264_),
    .B(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__mux2_1 _11188_ (.A0(\_152_[1] ),
    .A1(_05270_),
    .S(_01362_),
    .X(_05271_));
 sky130_fd_sc_hd__clkbuf_1 _11189_ (.A(_05271_),
    .X(_00724_));
 sky130_fd_sc_hd__nand2_1 _11190_ (.A(\_149_[1] ),
    .B(\_132_[1] ),
    .Y(_05272_));
 sky130_fd_sc_hd__o21a_1 _11191_ (.A1(_05264_),
    .A2(_05268_),
    .B1(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__nor2_1 _11192_ (.A(\_149_[2] ),
    .B(\_132_[2] ),
    .Y(_05274_));
 sky130_fd_sc_hd__nand2_1 _11193_ (.A(\_149_[2] ),
    .B(\_132_[2] ),
    .Y(_05275_));
 sky130_fd_sc_hd__and2b_1 _11194_ (.A_N(_05274_),
    .B(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__xnor2_1 _11195_ (.A(_05273_),
    .B(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__mux2_1 _11196_ (.A0(\_152_[2] ),
    .A1(_05277_),
    .S(_01362_),
    .X(_05278_));
 sky130_fd_sc_hd__clkbuf_1 _11197_ (.A(_05278_),
    .X(_00725_));
 sky130_fd_sc_hd__buf_4 _11198_ (.A(_05263_),
    .X(_05279_));
 sky130_fd_sc_hd__nor2_1 _11199_ (.A(\_149_[3] ),
    .B(\_132_[3] ),
    .Y(_05280_));
 sky130_fd_sc_hd__nand2_1 _11200_ (.A(\_149_[3] ),
    .B(\_132_[3] ),
    .Y(_05281_));
 sky130_fd_sc_hd__or2b_1 _11201_ (.A(_05280_),
    .B_N(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__o211a_1 _11202_ (.A1(_05264_),
    .A2(_05268_),
    .B1(_05275_),
    .C1(_05272_),
    .X(_05283_));
 sky130_fd_sc_hd__or3_1 _11203_ (.A(_05274_),
    .B(_05282_),
    .C(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__o21ai_1 _11204_ (.A1(_05274_),
    .A2(_05283_),
    .B1(_05282_),
    .Y(_05285_));
 sky130_fd_sc_hd__and2_1 _11205_ (.A(\_152_[3] ),
    .B(_01368_),
    .X(_05286_));
 sky130_fd_sc_hd__a31o_1 _11206_ (.A1(_05279_),
    .A2(_05284_),
    .A3(_05285_),
    .B1(_05286_),
    .X(_00726_));
 sky130_fd_sc_hd__or2_1 _11207_ (.A(\_149_[4] ),
    .B(\_132_[4] ),
    .X(_05287_));
 sky130_fd_sc_hd__nand2_1 _11208_ (.A(\_149_[4] ),
    .B(\_132_[4] ),
    .Y(_05288_));
 sky130_fd_sc_hd__nand2_1 _11209_ (.A(_05287_),
    .B(_05288_),
    .Y(_05289_));
 sky130_fd_sc_hd__o31a_1 _11210_ (.A1(_05274_),
    .A2(_05280_),
    .A3(_05283_),
    .B1(_05281_),
    .X(_05290_));
 sky130_fd_sc_hd__xor2_1 _11211_ (.A(_05289_),
    .B(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__mux2_1 _11212_ (.A0(\_152_[4] ),
    .A1(_05291_),
    .S(_01362_),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_1 _11213_ (.A(_05292_),
    .X(_00727_));
 sky130_fd_sc_hd__or2_1 _11214_ (.A(\_149_[5] ),
    .B(\_132_[5] ),
    .X(_05293_));
 sky130_fd_sc_hd__nand2_1 _11215_ (.A(\_149_[5] ),
    .B(\_132_[5] ),
    .Y(_05294_));
 sky130_fd_sc_hd__nand2_1 _11216_ (.A(_05293_),
    .B(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__o21ai_1 _11217_ (.A1(_05289_),
    .A2(_05290_),
    .B1(_05288_),
    .Y(_05296_));
 sky130_fd_sc_hd__xnor2_1 _11218_ (.A(_05295_),
    .B(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__mux2_1 _11219_ (.A0(\_152_[5] ),
    .A1(_05297_),
    .S(_01362_),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_1 _11220_ (.A(_05298_),
    .X(_00728_));
 sky130_fd_sc_hd__or2_1 _11221_ (.A(\_149_[6] ),
    .B(\_132_[6] ),
    .X(_05299_));
 sky130_fd_sc_hd__nand2_1 _11222_ (.A(\_149_[6] ),
    .B(\_132_[6] ),
    .Y(_05300_));
 sky130_fd_sc_hd__nand2_1 _11223_ (.A(_05299_),
    .B(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__nand3_1 _11224_ (.A(\_149_[4] ),
    .B(\_132_[4] ),
    .C(_05293_),
    .Y(_05302_));
 sky130_fd_sc_hd__o311a_1 _11225_ (.A1(_05289_),
    .A2(_05290_),
    .A3(_05295_),
    .B1(_05302_),
    .C1(_05294_),
    .X(_05303_));
 sky130_fd_sc_hd__xor2_1 _11226_ (.A(_05301_),
    .B(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__mux2_1 _11227_ (.A0(\_152_[6] ),
    .A1(_05304_),
    .S(_01362_),
    .X(_05305_));
 sky130_fd_sc_hd__clkbuf_1 _11228_ (.A(_05305_),
    .X(_00729_));
 sky130_fd_sc_hd__or2_1 _11229_ (.A(\_149_[7] ),
    .B(\_132_[7] ),
    .X(_05306_));
 sky130_fd_sc_hd__nand2_1 _11230_ (.A(\_149_[7] ),
    .B(\_132_[7] ),
    .Y(_05307_));
 sky130_fd_sc_hd__nand2_1 _11231_ (.A(_05306_),
    .B(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__o21ai_1 _11232_ (.A1(_05301_),
    .A2(_05303_),
    .B1(_05300_),
    .Y(_05309_));
 sky130_fd_sc_hd__xnor2_1 _11233_ (.A(_05308_),
    .B(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__mux2_1 _11234_ (.A0(\_152_[7] ),
    .A1(_05310_),
    .S(_01362_),
    .X(_05311_));
 sky130_fd_sc_hd__clkbuf_1 _11235_ (.A(_05311_),
    .X(_00730_));
 sky130_fd_sc_hd__or2_1 _11236_ (.A(\_149_[8] ),
    .B(\_132_[8] ),
    .X(_05312_));
 sky130_fd_sc_hd__nand2_1 _11237_ (.A(\_149_[8] ),
    .B(\_132_[8] ),
    .Y(_05313_));
 sky130_fd_sc_hd__nand2_1 _11238_ (.A(_05312_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__nand3_1 _11239_ (.A(\_149_[6] ),
    .B(\_132_[6] ),
    .C(_05306_),
    .Y(_05315_));
 sky130_fd_sc_hd__o311a_1 _11240_ (.A1(_05301_),
    .A2(_05303_),
    .A3(_05308_),
    .B1(_05315_),
    .C1(_05307_),
    .X(_05316_));
 sky130_fd_sc_hd__xor2_1 _11241_ (.A(_05314_),
    .B(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__buf_4 _11242_ (.A(_01361_),
    .X(_05318_));
 sky130_fd_sc_hd__mux2_1 _11243_ (.A0(\_152_[8] ),
    .A1(_05317_),
    .S(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__clkbuf_1 _11244_ (.A(_05319_),
    .X(_00731_));
 sky130_fd_sc_hd__nor2_1 _11245_ (.A(\_149_[9] ),
    .B(\_132_[9] ),
    .Y(_05320_));
 sky130_fd_sc_hd__nand2_1 _11246_ (.A(\_149_[9] ),
    .B(\_132_[9] ),
    .Y(_05321_));
 sky130_fd_sc_hd__or2b_1 _11247_ (.A(_05320_),
    .B_N(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__or2_1 _11248_ (.A(_05314_),
    .B(_05316_),
    .X(_05323_));
 sky130_fd_sc_hd__nand2_1 _11249_ (.A(_05313_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__xnor2_1 _11250_ (.A(_05322_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__mux2_1 _11251_ (.A0(\_152_[9] ),
    .A1(_05325_),
    .S(_05318_),
    .X(_05326_));
 sky130_fd_sc_hd__clkbuf_1 _11252_ (.A(_05326_),
    .X(_00732_));
 sky130_fd_sc_hd__or2_1 _11253_ (.A(\_149_[10] ),
    .B(\_132_[10] ),
    .X(_05327_));
 sky130_fd_sc_hd__nand2_1 _11254_ (.A(\_149_[10] ),
    .B(\_132_[10] ),
    .Y(_05328_));
 sky130_fd_sc_hd__and2_1 _11255_ (.A(_05327_),
    .B(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__inv_2 _11256_ (.A(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__a311o_2 _11257_ (.A1(_05313_),
    .A2(_05323_),
    .A3(_05321_),
    .B1(_05330_),
    .C1(_05320_),
    .X(_05331_));
 sky130_fd_sc_hd__a31o_1 _11258_ (.A1(_05313_),
    .A2(_05323_),
    .A3(_05321_),
    .B1(_05320_),
    .X(_05332_));
 sky130_fd_sc_hd__nand2_1 _11259_ (.A(_05330_),
    .B(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__and2_1 _11260_ (.A(\_152_[10] ),
    .B(_01368_),
    .X(_05334_));
 sky130_fd_sc_hd__a31o_1 _11261_ (.A1(_05279_),
    .A2(_05331_),
    .A3(_05333_),
    .B1(_05334_),
    .X(_00733_));
 sky130_fd_sc_hd__nor2_1 _11262_ (.A(\_149_[11] ),
    .B(\_132_[11] ),
    .Y(_05335_));
 sky130_fd_sc_hd__nand2_1 _11263_ (.A(\_149_[11] ),
    .B(\_132_[11] ),
    .Y(_05336_));
 sky130_fd_sc_hd__or2b_1 _11264_ (.A(_05335_),
    .B_N(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__nand2_1 _11265_ (.A(_05328_),
    .B(_05331_),
    .Y(_05338_));
 sky130_fd_sc_hd__xnor2_1 _11266_ (.A(_05337_),
    .B(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__mux2_1 _11267_ (.A0(\_152_[11] ),
    .A1(_05339_),
    .S(_05318_),
    .X(_05340_));
 sky130_fd_sc_hd__clkbuf_1 _11268_ (.A(_05340_),
    .X(_00734_));
 sky130_fd_sc_hd__or2_1 _11269_ (.A(\_149_[12] ),
    .B(\_132_[12] ),
    .X(_05341_));
 sky130_fd_sc_hd__nand2_1 _11270_ (.A(\_149_[12] ),
    .B(\_132_[12] ),
    .Y(_05342_));
 sky130_fd_sc_hd__nand2_1 _11271_ (.A(_05341_),
    .B(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__a311o_2 _11272_ (.A1(_05328_),
    .A2(_05331_),
    .A3(_05336_),
    .B1(_05343_),
    .C1(_05335_),
    .X(_05344_));
 sky130_fd_sc_hd__a31o_1 _11273_ (.A1(_05328_),
    .A2(_05331_),
    .A3(_05336_),
    .B1(_05335_),
    .X(_05345_));
 sky130_fd_sc_hd__nand2_1 _11274_ (.A(_05343_),
    .B(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__and2_1 _11275_ (.A(\_152_[12] ),
    .B(_01368_),
    .X(_05347_));
 sky130_fd_sc_hd__a31o_1 _11276_ (.A1(_05279_),
    .A2(_05344_),
    .A3(_05346_),
    .B1(_05347_),
    .X(_00735_));
 sky130_fd_sc_hd__nor2_1 _11277_ (.A(\_149_[13] ),
    .B(\_132_[13] ),
    .Y(_05348_));
 sky130_fd_sc_hd__nand2_1 _11278_ (.A(\_149_[13] ),
    .B(\_132_[13] ),
    .Y(_05349_));
 sky130_fd_sc_hd__or2b_1 _11279_ (.A(_05348_),
    .B_N(_05349_),
    .X(_05350_));
 sky130_fd_sc_hd__a21oi_1 _11280_ (.A1(_05342_),
    .A2(_05344_),
    .B1(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__buf_4 _11281_ (.A(_01367_),
    .X(_05352_));
 sky130_fd_sc_hd__a31o_1 _11282_ (.A1(_05342_),
    .A2(_05344_),
    .A3(_05350_),
    .B1(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__a2bb2o_1 _11283_ (.A1_N(_05351_),
    .A2_N(_05353_),
    .B1(\_152_[13] ),
    .B2(_05262_),
    .X(_00736_));
 sky130_fd_sc_hd__or2_1 _11284_ (.A(\_149_[14] ),
    .B(\_132_[14] ),
    .X(_05354_));
 sky130_fd_sc_hd__nand2_1 _11285_ (.A(\_149_[14] ),
    .B(\_132_[14] ),
    .Y(_05355_));
 sky130_fd_sc_hd__and2_1 _11286_ (.A(_05354_),
    .B(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__a31o_1 _11287_ (.A1(_05342_),
    .A2(_05344_),
    .A3(_05349_),
    .B1(_05348_),
    .X(_05357_));
 sky130_fd_sc_hd__xnor2_1 _11288_ (.A(_05356_),
    .B(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__mux2_1 _11289_ (.A0(\_152_[14] ),
    .A1(_05358_),
    .S(_05318_),
    .X(_05359_));
 sky130_fd_sc_hd__clkbuf_1 _11290_ (.A(_05359_),
    .X(_00737_));
 sky130_fd_sc_hd__nor2_1 _11291_ (.A(\_149_[15] ),
    .B(\_132_[15] ),
    .Y(_05360_));
 sky130_fd_sc_hd__nand2_1 _11292_ (.A(\_149_[15] ),
    .B(\_132_[15] ),
    .Y(_05361_));
 sky130_fd_sc_hd__or2b_1 _11293_ (.A(_05360_),
    .B_N(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__inv_2 _11294_ (.A(_05356_),
    .Y(_05363_));
 sky130_fd_sc_hd__a311o_1 _11295_ (.A1(_05342_),
    .A2(_05344_),
    .A3(_05349_),
    .B1(_05363_),
    .C1(_05348_),
    .X(_05364_));
 sky130_fd_sc_hd__nand2_1 _11296_ (.A(_05355_),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__xnor2_1 _11297_ (.A(_05362_),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__mux2_1 _11298_ (.A0(\_152_[15] ),
    .A1(_05366_),
    .S(_05318_),
    .X(_05367_));
 sky130_fd_sc_hd__clkbuf_1 _11299_ (.A(_05367_),
    .X(_00738_));
 sky130_fd_sc_hd__nand2_1 _11300_ (.A(\_149_[16] ),
    .B(\_132_[16] ),
    .Y(_05368_));
 sky130_fd_sc_hd__or2_1 _11301_ (.A(\_149_[16] ),
    .B(\_132_[16] ),
    .X(_05369_));
 sky130_fd_sc_hd__nand2_1 _11302_ (.A(_05368_),
    .B(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__a31o_1 _11303_ (.A1(_05355_),
    .A2(_05364_),
    .A3(_05361_),
    .B1(_05360_),
    .X(_05371_));
 sky130_fd_sc_hd__nand2_1 _11304_ (.A(_05370_),
    .B(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__a311o_1 _11305_ (.A1(_05355_),
    .A2(_05364_),
    .A3(_05361_),
    .B1(_05370_),
    .C1(_05360_),
    .X(_05373_));
 sky130_fd_sc_hd__and2_1 _11306_ (.A(\_152_[16] ),
    .B(_01368_),
    .X(_05374_));
 sky130_fd_sc_hd__a31o_1 _11307_ (.A1(_05279_),
    .A2(_05372_),
    .A3(_05373_),
    .B1(_05374_),
    .X(_00739_));
 sky130_fd_sc_hd__nor2_1 _11308_ (.A(\_149_[17] ),
    .B(\_132_[17] ),
    .Y(_05375_));
 sky130_fd_sc_hd__nand2_1 _11309_ (.A(\_149_[17] ),
    .B(\_132_[17] ),
    .Y(_05376_));
 sky130_fd_sc_hd__or2b_1 _11310_ (.A(_05375_),
    .B_N(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__nand2_1 _11311_ (.A(_05368_),
    .B(_05373_),
    .Y(_05378_));
 sky130_fd_sc_hd__xnor2_1 _11312_ (.A(_05377_),
    .B(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__mux2_1 _11313_ (.A0(\_152_[17] ),
    .A1(_05379_),
    .S(_05318_),
    .X(_05380_));
 sky130_fd_sc_hd__clkbuf_1 _11314_ (.A(_05380_),
    .X(_00740_));
 sky130_fd_sc_hd__nand2_1 _11315_ (.A(\_149_[18] ),
    .B(\_132_[18] ),
    .Y(_05381_));
 sky130_fd_sc_hd__or2_1 _11316_ (.A(\_149_[18] ),
    .B(\_132_[18] ),
    .X(_05382_));
 sky130_fd_sc_hd__nand2_1 _11317_ (.A(_05381_),
    .B(_05382_),
    .Y(_05383_));
 sky130_fd_sc_hd__a31o_1 _11318_ (.A1(_05368_),
    .A2(_05373_),
    .A3(_05376_),
    .B1(_05375_),
    .X(_05384_));
 sky130_fd_sc_hd__nand2_1 _11319_ (.A(_05383_),
    .B(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__a311o_1 _11320_ (.A1(_05368_),
    .A2(_05373_),
    .A3(_05376_),
    .B1(_05383_),
    .C1(_05375_),
    .X(_05386_));
 sky130_fd_sc_hd__and2_1 _11321_ (.A(\_152_[18] ),
    .B(_01368_),
    .X(_05387_));
 sky130_fd_sc_hd__a31o_1 _11322_ (.A1(_05279_),
    .A2(_05385_),
    .A3(_05386_),
    .B1(_05387_),
    .X(_00741_));
 sky130_fd_sc_hd__nor2_1 _11323_ (.A(\_149_[19] ),
    .B(\_132_[19] ),
    .Y(_05388_));
 sky130_fd_sc_hd__nand2_1 _11324_ (.A(\_149_[19] ),
    .B(\_132_[19] ),
    .Y(_05389_));
 sky130_fd_sc_hd__or2b_1 _11325_ (.A(_05388_),
    .B_N(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__nand2_1 _11326_ (.A(_05381_),
    .B(_05386_),
    .Y(_05391_));
 sky130_fd_sc_hd__xnor2_1 _11327_ (.A(_05390_),
    .B(_05391_),
    .Y(_05392_));
 sky130_fd_sc_hd__mux2_1 _11328_ (.A0(\_152_[19] ),
    .A1(_05392_),
    .S(_05318_),
    .X(_05393_));
 sky130_fd_sc_hd__clkbuf_1 _11329_ (.A(_05393_),
    .X(_00742_));
 sky130_fd_sc_hd__or2_1 _11330_ (.A(\_149_[20] ),
    .B(\_132_[20] ),
    .X(_05394_));
 sky130_fd_sc_hd__nand2_2 _11331_ (.A(\_149_[20] ),
    .B(\_132_[20] ),
    .Y(_05395_));
 sky130_fd_sc_hd__and2_1 _11332_ (.A(_05394_),
    .B(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__inv_2 _11333_ (.A(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__a31o_1 _11334_ (.A1(_05381_),
    .A2(_05386_),
    .A3(_05389_),
    .B1(_05388_),
    .X(_05398_));
 sky130_fd_sc_hd__nand2_1 _11335_ (.A(_05397_),
    .B(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__a311o_2 _11336_ (.A1(_05381_),
    .A2(_05386_),
    .A3(_05389_),
    .B1(_05397_),
    .C1(_05388_),
    .X(_05400_));
 sky130_fd_sc_hd__and2_1 _11337_ (.A(\_152_[20] ),
    .B(_01368_),
    .X(_05401_));
 sky130_fd_sc_hd__a31o_1 _11338_ (.A1(_05279_),
    .A2(_05399_),
    .A3(_05400_),
    .B1(_05401_),
    .X(_00743_));
 sky130_fd_sc_hd__nor2_1 _11339_ (.A(\_149_[21] ),
    .B(\_132_[21] ),
    .Y(_05402_));
 sky130_fd_sc_hd__nand2_1 _11340_ (.A(\_149_[21] ),
    .B(\_132_[21] ),
    .Y(_05403_));
 sky130_fd_sc_hd__or2b_1 _11341_ (.A(_05402_),
    .B_N(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__nand2_1 _11342_ (.A(_05395_),
    .B(_05400_),
    .Y(_05405_));
 sky130_fd_sc_hd__xnor2_1 _11343_ (.A(_05404_),
    .B(_05405_),
    .Y(_05406_));
 sky130_fd_sc_hd__mux2_1 _11344_ (.A0(\_152_[21] ),
    .A1(_05406_),
    .S(_05318_),
    .X(_05407_));
 sky130_fd_sc_hd__clkbuf_1 _11345_ (.A(_05407_),
    .X(_00744_));
 sky130_fd_sc_hd__nor2_1 _11346_ (.A(\_149_[22] ),
    .B(\_132_[22] ),
    .Y(_05408_));
 sky130_fd_sc_hd__and2_1 _11347_ (.A(\_149_[22] ),
    .B(\_132_[22] ),
    .X(_05409_));
 sky130_fd_sc_hd__nor2_1 _11348_ (.A(_05408_),
    .B(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__inv_2 _11349_ (.A(_05410_),
    .Y(_05411_));
 sky130_fd_sc_hd__a31o_1 _11350_ (.A1(_05395_),
    .A2(_05400_),
    .A3(_05403_),
    .B1(_05402_),
    .X(_05412_));
 sky130_fd_sc_hd__nand2_1 _11351_ (.A(_05411_),
    .B(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__a311oi_4 _11352_ (.A1(_05395_),
    .A2(_05400_),
    .A3(_05403_),
    .B1(_05411_),
    .C1(_05402_),
    .Y(_05414_));
 sky130_fd_sc_hd__nor2_1 _11353_ (.A(_05352_),
    .B(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__a22o_1 _11354_ (.A1(\_152_[22] ),
    .A2(_05262_),
    .B1(_05413_),
    .B2(_05415_),
    .X(_00745_));
 sky130_fd_sc_hd__or2_1 _11355_ (.A(\_149_[23] ),
    .B(\_132_[23] ),
    .X(_05416_));
 sky130_fd_sc_hd__nand2_1 _11356_ (.A(\_149_[23] ),
    .B(\_132_[23] ),
    .Y(_05417_));
 sky130_fd_sc_hd__o211a_1 _11357_ (.A1(_05409_),
    .A2(_05414_),
    .B1(_05416_),
    .C1(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__a211o_1 _11358_ (.A1(_05416_),
    .A2(_05417_),
    .B1(_05409_),
    .C1(_05414_),
    .X(_05419_));
 sky130_fd_sc_hd__nand2_1 _11359_ (.A(_05263_),
    .B(_05419_),
    .Y(_05420_));
 sky130_fd_sc_hd__a2bb2o_1 _11360_ (.A1_N(_05418_),
    .A2_N(_05420_),
    .B1(\_152_[23] ),
    .B2(_05262_),
    .X(_00746_));
 sky130_fd_sc_hd__xnor2_1 _11361_ (.A(\_149_[24] ),
    .B(\_132_[24] ),
    .Y(_05421_));
 sky130_fd_sc_hd__and2_1 _11362_ (.A(\_149_[23] ),
    .B(\_132_[23] ),
    .X(_05422_));
 sky130_fd_sc_hd__o31a_1 _11363_ (.A1(_05409_),
    .A2(_05414_),
    .A3(_05422_),
    .B1(_05416_),
    .X(_05423_));
 sky130_fd_sc_hd__xnor2_1 _11364_ (.A(_05421_),
    .B(_05423_),
    .Y(_05424_));
 sky130_fd_sc_hd__mux2_1 _11365_ (.A0(\_152_[24] ),
    .A1(_05424_),
    .S(_05318_),
    .X(_05425_));
 sky130_fd_sc_hd__clkbuf_1 _11366_ (.A(_05425_),
    .X(_00747_));
 sky130_fd_sc_hd__nand2_1 _11367_ (.A(\_149_[25] ),
    .B(\_132_[25] ),
    .Y(_05426_));
 sky130_fd_sc_hd__or2_1 _11368_ (.A(\_149_[25] ),
    .B(\_132_[25] ),
    .X(_05427_));
 sky130_fd_sc_hd__nand2_1 _11369_ (.A(_05426_),
    .B(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__and2b_1 _11370_ (.A_N(_05421_),
    .B(_05423_),
    .X(_05429_));
 sky130_fd_sc_hd__a21o_1 _11371_ (.A1(\_149_[24] ),
    .A2(\_132_[24] ),
    .B1(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__xnor2_1 _11372_ (.A(_05428_),
    .B(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__mux2_1 _11373_ (.A0(\_152_[25] ),
    .A1(_05431_),
    .S(_05318_),
    .X(_05432_));
 sky130_fd_sc_hd__clkbuf_1 _11374_ (.A(_05432_),
    .X(_00748_));
 sky130_fd_sc_hd__nor2_1 _11375_ (.A(\_149_[26] ),
    .B(\_132_[26] ),
    .Y(_05433_));
 sky130_fd_sc_hd__and2_1 _11376_ (.A(\_149_[26] ),
    .B(\_132_[26] ),
    .X(_05434_));
 sky130_fd_sc_hd__or2_1 _11377_ (.A(_05433_),
    .B(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__a22o_1 _11378_ (.A1(\_149_[24] ),
    .A2(\_132_[24] ),
    .B1(\_149_[25] ),
    .B2(\_132_[25] ),
    .X(_05436_));
 sky130_fd_sc_hd__o21a_1 _11379_ (.A1(_05429_),
    .A2(_05436_),
    .B1(_05427_),
    .X(_05437_));
 sky130_fd_sc_hd__xnor2_1 _11380_ (.A(_05435_),
    .B(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hd__clkbuf_4 _11381_ (.A(_01361_),
    .X(_05439_));
 sky130_fd_sc_hd__mux2_1 _11382_ (.A0(\_152_[26] ),
    .A1(_05438_),
    .S(_05439_),
    .X(_05440_));
 sky130_fd_sc_hd__clkbuf_1 _11383_ (.A(_05440_),
    .X(_00749_));
 sky130_fd_sc_hd__inv_2 _11384_ (.A(_05435_),
    .Y(_05441_));
 sky130_fd_sc_hd__and2_1 _11385_ (.A(_05441_),
    .B(_05437_),
    .X(_05442_));
 sky130_fd_sc_hd__nor2_1 _11386_ (.A(\_149_[27] ),
    .B(\_132_[27] ),
    .Y(_05443_));
 sky130_fd_sc_hd__and2_1 _11387_ (.A(\_149_[27] ),
    .B(\_132_[27] ),
    .X(_05444_));
 sky130_fd_sc_hd__nor2_1 _11388_ (.A(_05443_),
    .B(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__o21ai_1 _11389_ (.A1(_05434_),
    .A2(_05442_),
    .B1(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__o31a_1 _11390_ (.A1(_05434_),
    .A2(_05442_),
    .A3(_05445_),
    .B1(_05263_),
    .X(_05447_));
 sky130_fd_sc_hd__a22o_1 _11391_ (.A1(\_152_[27] ),
    .A2(_05262_),
    .B1(_05446_),
    .B2(_05447_),
    .X(_00750_));
 sky130_fd_sc_hd__and4bb_1 _11392_ (.A_N(_05421_),
    .B_N(_05428_),
    .C(_05441_),
    .D(_05445_),
    .X(_05448_));
 sky130_fd_sc_hd__o311a_1 _11393_ (.A1(_05409_),
    .A2(_05414_),
    .A3(_05422_),
    .B1(_05448_),
    .C1(_05416_),
    .X(_05449_));
 sky130_fd_sc_hd__and4_1 _11394_ (.A(_05427_),
    .B(_05441_),
    .C(_05436_),
    .D(_05445_),
    .X(_05450_));
 sky130_fd_sc_hd__and2b_1 _11395_ (.A_N(_05443_),
    .B(_05434_),
    .X(_05451_));
 sky130_fd_sc_hd__or4_1 _11396_ (.A(_05444_),
    .B(_05449_),
    .C(_05450_),
    .D(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__nand2_1 _11397_ (.A(\_149_[28] ),
    .B(\_132_[28] ),
    .Y(_05453_));
 sky130_fd_sc_hd__or2_1 _11398_ (.A(\_149_[28] ),
    .B(\_132_[28] ),
    .X(_05454_));
 sky130_fd_sc_hd__nand2_1 _11399_ (.A(_05453_),
    .B(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__xnor2_1 _11400_ (.A(_05452_),
    .B(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__mux2_1 _11401_ (.A0(\_152_[28] ),
    .A1(_05456_),
    .S(_05439_),
    .X(_05457_));
 sky130_fd_sc_hd__clkbuf_1 _11402_ (.A(_05457_),
    .X(_00751_));
 sky130_fd_sc_hd__nand2_1 _11403_ (.A(\_149_[29] ),
    .B(\_132_[29] ),
    .Y(_05458_));
 sky130_fd_sc_hd__or2_1 _11404_ (.A(\_149_[29] ),
    .B(\_132_[29] ),
    .X(_05459_));
 sky130_fd_sc_hd__a21boi_1 _11405_ (.A1(_05452_),
    .A2(_05454_),
    .B1_N(_05453_),
    .Y(_05460_));
 sky130_fd_sc_hd__and3_1 _11406_ (.A(_05458_),
    .B(_05459_),
    .C(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__a21o_1 _11407_ (.A1(_05458_),
    .A2(_05459_),
    .B1(_05460_),
    .X(_05462_));
 sky130_fd_sc_hd__nand2_1 _11408_ (.A(_05263_),
    .B(_05462_),
    .Y(_05463_));
 sky130_fd_sc_hd__o22a_1 _11409_ (.A1(\_152_[29] ),
    .A2(_05279_),
    .B1(_05461_),
    .B2(_05463_),
    .X(_00752_));
 sky130_fd_sc_hd__and2_1 _11410_ (.A(\_149_[30] ),
    .B(\_132_[30] ),
    .X(_05464_));
 sky130_fd_sc_hd__or2_1 _11411_ (.A(\_149_[30] ),
    .B(\_132_[30] ),
    .X(_05465_));
 sky130_fd_sc_hd__or2b_1 _11412_ (.A(_05464_),
    .B_N(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__nor2_1 _11413_ (.A(\_149_[29] ),
    .B(\_132_[29] ),
    .Y(_05467_));
 sky130_fd_sc_hd__o21ai_1 _11414_ (.A1(_05467_),
    .A2(_05460_),
    .B1(_05458_),
    .Y(_05468_));
 sky130_fd_sc_hd__xnor2_1 _11415_ (.A(_05466_),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__mux2_1 _11416_ (.A0(\_152_[30] ),
    .A1(_05469_),
    .S(_05439_),
    .X(_05470_));
 sky130_fd_sc_hd__clkbuf_1 _11417_ (.A(_05470_),
    .X(_00753_));
 sky130_fd_sc_hd__a21o_1 _11418_ (.A1(_05465_),
    .A2(_05468_),
    .B1(_05464_),
    .X(_05471_));
 sky130_fd_sc_hd__xnor2_1 _11419_ (.A(\_149_[31] ),
    .B(\_132_[31] ),
    .Y(_05472_));
 sky130_fd_sc_hd__xnor2_1 _11420_ (.A(_05471_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__mux2_1 _11421_ (.A0(\_152_[31] ),
    .A1(_05473_),
    .S(_05439_),
    .X(_05474_));
 sky130_fd_sc_hd__clkbuf_1 _11422_ (.A(_05474_),
    .X(_00754_));
 sky130_fd_sc_hd__xnor2_1 _11423_ (.A(\_118_[7] ),
    .B(\_118_[3] ),
    .Y(_05475_));
 sky130_fd_sc_hd__xnor2_1 _11424_ (.A(\_118_[18] ),
    .B(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_1 _11425_ (.A(\_116_[0] ),
    .B(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__o21a_1 _11426_ (.A1(\_116_[0] ),
    .A2(_05476_),
    .B1(_05263_),
    .X(_05478_));
 sky130_fd_sc_hd__a22o_1 _11427_ (.A1(\_149_[0] ),
    .A2(_05352_),
    .B1(_05477_),
    .B2(_05478_),
    .X(_00755_));
 sky130_fd_sc_hd__xnor2_1 _11428_ (.A(\_118_[8] ),
    .B(\_118_[4] ),
    .Y(_05479_));
 sky130_fd_sc_hd__xnor2_1 _11429_ (.A(\_118_[19] ),
    .B(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__xnor2_1 _11430_ (.A(\_116_[1] ),
    .B(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__xor2_1 _11431_ (.A(_05477_),
    .B(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__mux2_1 _11432_ (.A0(\_149_[1] ),
    .A1(_05482_),
    .S(_05439_),
    .X(_05483_));
 sky130_fd_sc_hd__clkbuf_1 _11433_ (.A(_05483_),
    .X(_00756_));
 sky130_fd_sc_hd__xnor2_1 _11434_ (.A(\_118_[9] ),
    .B(\_118_[5] ),
    .Y(_05484_));
 sky130_fd_sc_hd__xnor2_1 _11435_ (.A(\_118_[20] ),
    .B(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__and2_1 _11436_ (.A(\_116_[2] ),
    .B(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__or2_1 _11437_ (.A(\_116_[2] ),
    .B(_05485_),
    .X(_05487_));
 sky130_fd_sc_hd__or2b_1 _11438_ (.A(_05486_),
    .B_N(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__nand2_1 _11439_ (.A(\_116_[1] ),
    .B(_05480_),
    .Y(_05489_));
 sky130_fd_sc_hd__o21ai_1 _11440_ (.A1(_05477_),
    .A2(_05481_),
    .B1(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__xnor2_1 _11441_ (.A(_05488_),
    .B(_05490_),
    .Y(_05491_));
 sky130_fd_sc_hd__mux2_1 _11442_ (.A0(\_149_[2] ),
    .A1(_05491_),
    .S(_05439_),
    .X(_05492_));
 sky130_fd_sc_hd__clkbuf_1 _11443_ (.A(_05492_),
    .X(_00757_));
 sky130_fd_sc_hd__xnor2_1 _11444_ (.A(\_118_[10] ),
    .B(\_118_[6] ),
    .Y(_05493_));
 sky130_fd_sc_hd__xnor2_1 _11445_ (.A(\_118_[21] ),
    .B(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__and2_1 _11446_ (.A(\_116_[3] ),
    .B(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__or2_1 _11447_ (.A(\_116_[3] ),
    .B(_05494_),
    .X(_05496_));
 sky130_fd_sc_hd__or2b_1 _11448_ (.A(_05495_),
    .B_N(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__a21o_1 _11449_ (.A1(_05487_),
    .A2(_05490_),
    .B1(_05486_),
    .X(_05498_));
 sky130_fd_sc_hd__xnor2_1 _11450_ (.A(_05497_),
    .B(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__mux2_1 _11451_ (.A0(\_149_[3] ),
    .A1(_05499_),
    .S(_05439_),
    .X(_05500_));
 sky130_fd_sc_hd__clkbuf_1 _11452_ (.A(_05500_),
    .X(_00758_));
 sky130_fd_sc_hd__a21oi_2 _11453_ (.A1(_05496_),
    .A2(_05498_),
    .B1(_05495_),
    .Y(_05501_));
 sky130_fd_sc_hd__xnor2_1 _11454_ (.A(\_118_[22] ),
    .B(\_118_[11] ),
    .Y(_05502_));
 sky130_fd_sc_hd__xnor2_1 _11455_ (.A(\_118_[7] ),
    .B(_05502_),
    .Y(_05503_));
 sky130_fd_sc_hd__nand2_1 _11456_ (.A(\_116_[4] ),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__or2_1 _11457_ (.A(\_116_[4] ),
    .B(_05503_),
    .X(_05505_));
 sky130_fd_sc_hd__nand2_1 _11458_ (.A(_05504_),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__xor2_1 _11459_ (.A(_05501_),
    .B(_05506_),
    .X(_05507_));
 sky130_fd_sc_hd__mux2_1 _11460_ (.A0(\_149_[4] ),
    .A1(_05507_),
    .S(_05439_),
    .X(_05508_));
 sky130_fd_sc_hd__clkbuf_1 _11461_ (.A(_05508_),
    .X(_00759_));
 sky130_fd_sc_hd__xnor2_1 _11462_ (.A(\_118_[23] ),
    .B(\_118_[12] ),
    .Y(_05509_));
 sky130_fd_sc_hd__xnor2_1 _11463_ (.A(\_118_[8] ),
    .B(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__xnor2_1 _11464_ (.A(\_116_[5] ),
    .B(_05510_),
    .Y(_05511_));
 sky130_fd_sc_hd__o21ai_1 _11465_ (.A1(_05501_),
    .A2(_05506_),
    .B1(_05504_),
    .Y(_05512_));
 sky130_fd_sc_hd__xnor2_1 _11466_ (.A(_05511_),
    .B(_05512_),
    .Y(_05513_));
 sky130_fd_sc_hd__mux2_1 _11467_ (.A0(\_149_[5] ),
    .A1(_05513_),
    .S(_05439_),
    .X(_05514_));
 sky130_fd_sc_hd__clkbuf_1 _11468_ (.A(_05514_),
    .X(_00760_));
 sky130_fd_sc_hd__xnor2_1 _11469_ (.A(\_118_[24] ),
    .B(\_118_[13] ),
    .Y(_05515_));
 sky130_fd_sc_hd__xnor2_1 _11470_ (.A(\_118_[9] ),
    .B(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__nand2_1 _11471_ (.A(\_116_[6] ),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__or2_1 _11472_ (.A(\_116_[6] ),
    .B(_05516_),
    .X(_05518_));
 sky130_fd_sc_hd__nand2_1 _11473_ (.A(_05517_),
    .B(_05518_),
    .Y(_05519_));
 sky130_fd_sc_hd__or2_1 _11474_ (.A(_05506_),
    .B(_05511_),
    .X(_05520_));
 sky130_fd_sc_hd__a22o_1 _11475_ (.A1(\_116_[4] ),
    .A2(_05503_),
    .B1(_05510_),
    .B2(\_116_[5] ),
    .X(_05521_));
 sky130_fd_sc_hd__o21ai_1 _11476_ (.A1(\_116_[5] ),
    .A2(_05510_),
    .B1(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__o21ai_1 _11477_ (.A1(_05501_),
    .A2(_05520_),
    .B1(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__xnor2_1 _11478_ (.A(_05519_),
    .B(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__mux2_1 _11479_ (.A0(\_149_[6] ),
    .A1(_05524_),
    .S(_05439_),
    .X(_05525_));
 sky130_fd_sc_hd__clkbuf_1 _11480_ (.A(_05525_),
    .X(_00761_));
 sky130_fd_sc_hd__xnor2_1 _11481_ (.A(\_118_[25] ),
    .B(\_118_[14] ),
    .Y(_05526_));
 sky130_fd_sc_hd__xnor2_1 _11482_ (.A(\_118_[10] ),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__nor2_1 _11483_ (.A(\_116_[7] ),
    .B(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__nand2_1 _11484_ (.A(\_116_[7] ),
    .B(_05527_),
    .Y(_05529_));
 sky130_fd_sc_hd__or2b_1 _11485_ (.A(_05528_),
    .B_N(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__a21bo_1 _11486_ (.A1(_05518_),
    .A2(_05523_),
    .B1_N(_05517_),
    .X(_05531_));
 sky130_fd_sc_hd__xnor2_1 _11487_ (.A(_05530_),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__buf_4 _11488_ (.A(_01361_),
    .X(_05533_));
 sky130_fd_sc_hd__mux2_1 _11489_ (.A0(\_149_[7] ),
    .A1(_05532_),
    .S(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__clkbuf_1 _11490_ (.A(_05534_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _11491_ (.A(_05519_),
    .B(_05530_),
    .X(_05535_));
 sky130_fd_sc_hd__or2_1 _11492_ (.A(_05520_),
    .B(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__o21a_1 _11493_ (.A1(_05517_),
    .A2(_05528_),
    .B1(_05529_),
    .X(_05537_));
 sky130_fd_sc_hd__or2_1 _11494_ (.A(_05522_),
    .B(_05535_),
    .X(_05538_));
 sky130_fd_sc_hd__o211a_1 _11495_ (.A1(_05501_),
    .A2(_05536_),
    .B1(_05537_),
    .C1(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__xnor2_1 _11496_ (.A(\_118_[26] ),
    .B(\_118_[15] ),
    .Y(_05540_));
 sky130_fd_sc_hd__xnor2_1 _11497_ (.A(\_118_[11] ),
    .B(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hd__nand2_1 _11498_ (.A(\_116_[8] ),
    .B(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__or2_1 _11499_ (.A(\_116_[8] ),
    .B(_05541_),
    .X(_05543_));
 sky130_fd_sc_hd__nand2_1 _11500_ (.A(_05542_),
    .B(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__xor2_1 _11501_ (.A(_05539_),
    .B(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__mux2_1 _11502_ (.A0(\_149_[8] ),
    .A1(_05545_),
    .S(_05533_),
    .X(_05546_));
 sky130_fd_sc_hd__clkbuf_1 _11503_ (.A(_05546_),
    .X(_00763_));
 sky130_fd_sc_hd__xnor2_1 _11504_ (.A(\_118_[27] ),
    .B(\_118_[16] ),
    .Y(_05547_));
 sky130_fd_sc_hd__xnor2_1 _11505_ (.A(\_118_[12] ),
    .B(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__nand2_1 _11506_ (.A(\_116_[9] ),
    .B(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__nor2_1 _11507_ (.A(\_116_[9] ),
    .B(_05548_),
    .Y(_05550_));
 sky130_fd_sc_hd__inv_2 _11508_ (.A(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__nand2_1 _11509_ (.A(_05549_),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__o21ai_1 _11510_ (.A1(_05539_),
    .A2(_05544_),
    .B1(_05542_),
    .Y(_05553_));
 sky130_fd_sc_hd__xnor2_1 _11511_ (.A(_05552_),
    .B(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__mux2_1 _11512_ (.A0(\_149_[9] ),
    .A1(_05554_),
    .S(_05533_),
    .X(_05555_));
 sky130_fd_sc_hd__clkbuf_1 _11513_ (.A(_05555_),
    .X(_00764_));
 sky130_fd_sc_hd__xnor2_1 _11514_ (.A(\_118_[28] ),
    .B(\_118_[17] ),
    .Y(_05556_));
 sky130_fd_sc_hd__xnor2_1 _11515_ (.A(\_118_[13] ),
    .B(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__nand2_1 _11516_ (.A(\_116_[10] ),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__or2_1 _11517_ (.A(\_116_[10] ),
    .B(_05557_),
    .X(_05559_));
 sky130_fd_sc_hd__nand2_1 _11518_ (.A(_05558_),
    .B(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__a21o_1 _11519_ (.A1(_05542_),
    .A2(_05549_),
    .B1(_05550_),
    .X(_05561_));
 sky130_fd_sc_hd__o31a_1 _11520_ (.A1(_05539_),
    .A2(_05544_),
    .A3(_05552_),
    .B1(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__xor2_1 _11521_ (.A(_05560_),
    .B(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__mux2_1 _11522_ (.A0(\_149_[10] ),
    .A1(_05563_),
    .S(_05533_),
    .X(_05564_));
 sky130_fd_sc_hd__clkbuf_1 _11523_ (.A(_05564_),
    .X(_00765_));
 sky130_fd_sc_hd__xnor2_1 _11524_ (.A(\_118_[14] ),
    .B(\_118_[29] ),
    .Y(_05565_));
 sky130_fd_sc_hd__xnor2_1 _11525_ (.A(\_118_[18] ),
    .B(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__nand2_1 _11526_ (.A(\_116_[11] ),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__nor2_1 _11527_ (.A(\_116_[11] ),
    .B(_05566_),
    .Y(_05568_));
 sky130_fd_sc_hd__inv_2 _11528_ (.A(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__nand2_1 _11529_ (.A(_05567_),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__o21ai_1 _11530_ (.A1(_05560_),
    .A2(_05562_),
    .B1(_05558_),
    .Y(_05571_));
 sky130_fd_sc_hd__xnor2_1 _11531_ (.A(_05570_),
    .B(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__mux2_1 _11532_ (.A0(\_149_[11] ),
    .A1(_05572_),
    .S(_05533_),
    .X(_05573_));
 sky130_fd_sc_hd__clkbuf_1 _11533_ (.A(_05573_),
    .X(_00766_));
 sky130_fd_sc_hd__xnor2_1 _11534_ (.A(\_118_[15] ),
    .B(\_118_[30] ),
    .Y(_05574_));
 sky130_fd_sc_hd__xnor2_1 _11535_ (.A(\_118_[19] ),
    .B(_05574_),
    .Y(_05575_));
 sky130_fd_sc_hd__nand2_1 _11536_ (.A(\_116_[12] ),
    .B(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__or2_1 _11537_ (.A(\_116_[12] ),
    .B(_05575_),
    .X(_05577_));
 sky130_fd_sc_hd__nand2_1 _11538_ (.A(_05576_),
    .B(_05577_),
    .Y(_05578_));
 sky130_fd_sc_hd__a21o_1 _11539_ (.A1(_05558_),
    .A2(_05567_),
    .B1(_05568_),
    .X(_05579_));
 sky130_fd_sc_hd__o31a_1 _11540_ (.A1(_05560_),
    .A2(_05562_),
    .A3(_05570_),
    .B1(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__xor2_1 _11541_ (.A(_05578_),
    .B(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__mux2_1 _11542_ (.A0(\_149_[12] ),
    .A1(_05581_),
    .S(_05533_),
    .X(_05582_));
 sky130_fd_sc_hd__clkbuf_1 _11543_ (.A(_05582_),
    .X(_00767_));
 sky130_fd_sc_hd__xnor2_1 _11544_ (.A(\_118_[16] ),
    .B(\_118_[31] ),
    .Y(_05583_));
 sky130_fd_sc_hd__xnor2_1 _11545_ (.A(\_118_[20] ),
    .B(_05583_),
    .Y(_05584_));
 sky130_fd_sc_hd__nor2_1 _11546_ (.A(\_116_[13] ),
    .B(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__nand2_1 _11547_ (.A(\_116_[13] ),
    .B(_05584_),
    .Y(_05586_));
 sky130_fd_sc_hd__or2b_1 _11548_ (.A(_05585_),
    .B_N(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__o21ai_1 _11549_ (.A1(_05578_),
    .A2(_05580_),
    .B1(_05576_),
    .Y(_05588_));
 sky130_fd_sc_hd__xnor2_1 _11550_ (.A(_05587_),
    .B(_05588_),
    .Y(_05589_));
 sky130_fd_sc_hd__mux2_1 _11551_ (.A0(\_149_[13] ),
    .A1(_05589_),
    .S(_05533_),
    .X(_05590_));
 sky130_fd_sc_hd__clkbuf_1 _11552_ (.A(_05590_),
    .X(_00768_));
 sky130_fd_sc_hd__xnor2_1 _11553_ (.A(\_118_[17] ),
    .B(\_118_[0] ),
    .Y(_05591_));
 sky130_fd_sc_hd__xnor2_1 _11554_ (.A(\_118_[21] ),
    .B(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__nand2_1 _11555_ (.A(\_116_[14] ),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__or2_1 _11556_ (.A(\_116_[14] ),
    .B(_05592_),
    .X(_05594_));
 sky130_fd_sc_hd__nand2_1 _11557_ (.A(_05593_),
    .B(_05594_),
    .Y(_05595_));
 sky130_fd_sc_hd__a21o_1 _11558_ (.A1(_05576_),
    .A2(_05586_),
    .B1(_05585_),
    .X(_05596_));
 sky130_fd_sc_hd__o31a_1 _11559_ (.A1(_05578_),
    .A2(_05580_),
    .A3(_05587_),
    .B1(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__xor2_1 _11560_ (.A(_05595_),
    .B(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__mux2_1 _11561_ (.A0(\_149_[14] ),
    .A1(_05598_),
    .S(_05533_),
    .X(_05599_));
 sky130_fd_sc_hd__clkbuf_1 _11562_ (.A(_05599_),
    .X(_00769_));
 sky130_fd_sc_hd__xnor2_1 _11563_ (.A(\_118_[22] ),
    .B(\_118_[1] ),
    .Y(_05600_));
 sky130_fd_sc_hd__xnor2_1 _11564_ (.A(\_118_[18] ),
    .B(_05600_),
    .Y(_05601_));
 sky130_fd_sc_hd__nor2_1 _11565_ (.A(\_116_[15] ),
    .B(_05601_),
    .Y(_05602_));
 sky130_fd_sc_hd__nand2_1 _11566_ (.A(\_116_[15] ),
    .B(_05601_),
    .Y(_05603_));
 sky130_fd_sc_hd__or2b_1 _11567_ (.A(_05602_),
    .B_N(_05603_),
    .X(_05604_));
 sky130_fd_sc_hd__o21ai_1 _11568_ (.A1(_05595_),
    .A2(_05597_),
    .B1(_05593_),
    .Y(_05605_));
 sky130_fd_sc_hd__xnor2_1 _11569_ (.A(_05604_),
    .B(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__mux2_1 _11570_ (.A0(\_149_[15] ),
    .A1(_05606_),
    .S(_05533_),
    .X(_05607_));
 sky130_fd_sc_hd__clkbuf_1 _11571_ (.A(_05607_),
    .X(_00770_));
 sky130_fd_sc_hd__xnor2_1 _11572_ (.A(\_118_[23] ),
    .B(\_118_[2] ),
    .Y(_05608_));
 sky130_fd_sc_hd__xnor2_1 _11573_ (.A(\_118_[19] ),
    .B(_05608_),
    .Y(_05609_));
 sky130_fd_sc_hd__nand2_1 _11574_ (.A(\_116_[16] ),
    .B(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__or2_1 _11575_ (.A(\_116_[16] ),
    .B(_05609_),
    .X(_05611_));
 sky130_fd_sc_hd__nand2_1 _11576_ (.A(_05610_),
    .B(_05611_),
    .Y(_05612_));
 sky130_fd_sc_hd__a21o_1 _11577_ (.A1(_05593_),
    .A2(_05603_),
    .B1(_05602_),
    .X(_05613_));
 sky130_fd_sc_hd__o31a_1 _11578_ (.A1(_05595_),
    .A2(_05597_),
    .A3(_05604_),
    .B1(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__xor2_1 _11579_ (.A(_05612_),
    .B(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__mux2_1 _11580_ (.A0(\_149_[16] ),
    .A1(_05615_),
    .S(_05533_),
    .X(_05616_));
 sky130_fd_sc_hd__clkbuf_1 _11581_ (.A(_05616_),
    .X(_00771_));
 sky130_fd_sc_hd__xnor2_1 _11582_ (.A(\_118_[20] ),
    .B(\_118_[24] ),
    .Y(_05617_));
 sky130_fd_sc_hd__xnor2_1 _11583_ (.A(\_118_[3] ),
    .B(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand2_1 _11584_ (.A(\_116_[17] ),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__nor2_1 _11585_ (.A(\_116_[17] ),
    .B(_05618_),
    .Y(_05620_));
 sky130_fd_sc_hd__inv_2 _11586_ (.A(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__nand2_1 _11587_ (.A(_05619_),
    .B(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hd__o21ai_1 _11588_ (.A1(_05612_),
    .A2(_05614_),
    .B1(_05610_),
    .Y(_05623_));
 sky130_fd_sc_hd__xnor2_1 _11589_ (.A(_05622_),
    .B(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__buf_4 _11590_ (.A(_01361_),
    .X(_05625_));
 sky130_fd_sc_hd__mux2_1 _11591_ (.A0(\_149_[17] ),
    .A1(_05624_),
    .S(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__clkbuf_1 _11592_ (.A(_05626_),
    .X(_00772_));
 sky130_fd_sc_hd__xnor2_1 _11593_ (.A(\_118_[21] ),
    .B(\_118_[25] ),
    .Y(_05627_));
 sky130_fd_sc_hd__xnor2_1 _11594_ (.A(\_118_[4] ),
    .B(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__nand2_1 _11595_ (.A(\_116_[18] ),
    .B(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__or2_1 _11596_ (.A(\_116_[18] ),
    .B(_05628_),
    .X(_05630_));
 sky130_fd_sc_hd__nand2_1 _11597_ (.A(_05629_),
    .B(_05630_),
    .Y(_05631_));
 sky130_fd_sc_hd__a21o_1 _11598_ (.A1(_05610_),
    .A2(_05619_),
    .B1(_05620_),
    .X(_05632_));
 sky130_fd_sc_hd__o31a_1 _11599_ (.A1(_05612_),
    .A2(_05614_),
    .A3(_05622_),
    .B1(_05632_),
    .X(_05633_));
 sky130_fd_sc_hd__or2_1 _11600_ (.A(_05631_),
    .B(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__a21oi_1 _11601_ (.A1(_05631_),
    .A2(_05633_),
    .B1(_05352_),
    .Y(_05635_));
 sky130_fd_sc_hd__a22o_1 _11602_ (.A1(\_149_[18] ),
    .A2(_05352_),
    .B1(_05634_),
    .B2(_05635_),
    .X(_00773_));
 sky130_fd_sc_hd__xnor2_1 _11603_ (.A(\_118_[22] ),
    .B(\_118_[26] ),
    .Y(_05636_));
 sky130_fd_sc_hd__xnor2_1 _11604_ (.A(\_118_[5] ),
    .B(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_1 _11605_ (.A(\_116_[19] ),
    .B(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__nor2_1 _11606_ (.A(\_116_[19] ),
    .B(_05637_),
    .Y(_05639_));
 sky130_fd_sc_hd__inv_2 _11607_ (.A(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__nand2_1 _11608_ (.A(_05638_),
    .B(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__a21oi_1 _11609_ (.A1(_05629_),
    .A2(_05634_),
    .B1(_05641_),
    .Y(_05642_));
 sky130_fd_sc_hd__a31o_1 _11610_ (.A1(_05629_),
    .A2(_05634_),
    .A3(_05641_),
    .B1(_05352_),
    .X(_05643_));
 sky130_fd_sc_hd__a2bb2o_1 _11611_ (.A1_N(_05642_),
    .A2_N(_05643_),
    .B1(\_149_[19] ),
    .B2(_05262_),
    .X(_00774_));
 sky130_fd_sc_hd__xnor2_1 _11612_ (.A(\_118_[23] ),
    .B(\_118_[27] ),
    .Y(_05644_));
 sky130_fd_sc_hd__xnor2_1 _11613_ (.A(\_118_[6] ),
    .B(_05644_),
    .Y(_05645_));
 sky130_fd_sc_hd__nand2_1 _11614_ (.A(\_116_[20] ),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__or2_1 _11615_ (.A(\_116_[20] ),
    .B(_05645_),
    .X(_05647_));
 sky130_fd_sc_hd__nand2_1 _11616_ (.A(_05646_),
    .B(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__o211a_1 _11617_ (.A1(_05631_),
    .A2(_05633_),
    .B1(_05638_),
    .C1(_05629_),
    .X(_05649_));
 sky130_fd_sc_hd__or3_1 _11618_ (.A(_05639_),
    .B(_05648_),
    .C(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__o21ai_1 _11619_ (.A1(_05639_),
    .A2(_05649_),
    .B1(_05648_),
    .Y(_05651_));
 sky130_fd_sc_hd__and3_1 _11620_ (.A(_01362_),
    .B(_05650_),
    .C(_05651_),
    .X(_05652_));
 sky130_fd_sc_hd__a21o_1 _11621_ (.A1(\_149_[20] ),
    .A2(_05262_),
    .B1(_05652_),
    .X(_00775_));
 sky130_fd_sc_hd__xnor2_1 _11622_ (.A(\_118_[24] ),
    .B(\_118_[28] ),
    .Y(_05653_));
 sky130_fd_sc_hd__xnor2_1 _11623_ (.A(\_118_[7] ),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand2_1 _11624_ (.A(\_116_[21] ),
    .B(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__nor2_1 _11625_ (.A(\_116_[21] ),
    .B(_05654_),
    .Y(_05656_));
 sky130_fd_sc_hd__inv_2 _11626_ (.A(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__nand2_1 _11627_ (.A(_05655_),
    .B(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__a21oi_1 _11628_ (.A1(_05646_),
    .A2(_05650_),
    .B1(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__a31o_1 _11629_ (.A1(_05646_),
    .A2(_05650_),
    .A3(_05658_),
    .B1(_05352_),
    .X(_05660_));
 sky130_fd_sc_hd__a2bb2o_1 _11630_ (.A1_N(_05659_),
    .A2_N(_05660_),
    .B1(\_149_[21] ),
    .B2(_05262_),
    .X(_00776_));
 sky130_fd_sc_hd__xnor2_1 _11631_ (.A(\_118_[25] ),
    .B(\_118_[29] ),
    .Y(_05661_));
 sky130_fd_sc_hd__xnor2_1 _11632_ (.A(\_118_[8] ),
    .B(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__nand2_1 _11633_ (.A(\_116_[22] ),
    .B(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__or2_1 _11634_ (.A(\_116_[22] ),
    .B(_05662_),
    .X(_05664_));
 sky130_fd_sc_hd__nand2_1 _11635_ (.A(_05663_),
    .B(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__a21o_1 _11636_ (.A1(_05646_),
    .A2(_05655_),
    .B1(_05656_),
    .X(_05666_));
 sky130_fd_sc_hd__o41a_1 _11637_ (.A1(_05639_),
    .A2(_05648_),
    .A3(_05649_),
    .A4(_05658_),
    .B1(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__xor2_1 _11638_ (.A(_05665_),
    .B(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__mux2_1 _11639_ (.A0(\_149_[22] ),
    .A1(_05668_),
    .S(_05625_),
    .X(_05669_));
 sky130_fd_sc_hd__clkbuf_1 _11640_ (.A(_05669_),
    .X(_00777_));
 sky130_fd_sc_hd__xnor2_1 _11641_ (.A(\_118_[26] ),
    .B(\_118_[30] ),
    .Y(_05670_));
 sky130_fd_sc_hd__xnor2_1 _11642_ (.A(\_118_[9] ),
    .B(_05670_),
    .Y(_05671_));
 sky130_fd_sc_hd__xnor2_1 _11643_ (.A(\_116_[23] ),
    .B(_05671_),
    .Y(_05672_));
 sky130_fd_sc_hd__o21ai_1 _11644_ (.A1(_05665_),
    .A2(_05667_),
    .B1(_05663_),
    .Y(_05673_));
 sky130_fd_sc_hd__xnor2_1 _11645_ (.A(_05672_),
    .B(_05673_),
    .Y(_05674_));
 sky130_fd_sc_hd__mux2_1 _11646_ (.A0(\_149_[23] ),
    .A1(_05674_),
    .S(_05625_),
    .X(_05675_));
 sky130_fd_sc_hd__clkbuf_1 _11647_ (.A(_05675_),
    .X(_00778_));
 sky130_fd_sc_hd__xnor2_1 _11648_ (.A(\_118_[27] ),
    .B(\_118_[31] ),
    .Y(_05676_));
 sky130_fd_sc_hd__xnor2_1 _11649_ (.A(\_118_[10] ),
    .B(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__nand2_1 _11650_ (.A(\_116_[24] ),
    .B(_05677_),
    .Y(_05678_));
 sky130_fd_sc_hd__or2_1 _11651_ (.A(\_116_[24] ),
    .B(_05677_),
    .X(_05679_));
 sky130_fd_sc_hd__nand2_1 _11652_ (.A(_05678_),
    .B(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__a22o_1 _11653_ (.A1(\_116_[22] ),
    .A2(_05662_),
    .B1(_05671_),
    .B2(\_116_[23] ),
    .X(_05681_));
 sky130_fd_sc_hd__o21ai_1 _11654_ (.A1(\_116_[23] ),
    .A2(_05671_),
    .B1(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__o31a_1 _11655_ (.A1(_05665_),
    .A2(_05667_),
    .A3(_05672_),
    .B1(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__or2_1 _11656_ (.A(_05680_),
    .B(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__a21oi_1 _11657_ (.A1(_05680_),
    .A2(_05683_),
    .B1(_05352_),
    .Y(_05685_));
 sky130_fd_sc_hd__a22o_1 _11658_ (.A1(\_149_[24] ),
    .A2(_05352_),
    .B1(_05684_),
    .B2(_05685_),
    .X(_00779_));
 sky130_fd_sc_hd__xnor2_1 _11659_ (.A(\_118_[28] ),
    .B(\_118_[0] ),
    .Y(_05686_));
 sky130_fd_sc_hd__xnor2_2 _11660_ (.A(\_118_[11] ),
    .B(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__xnor2_1 _11661_ (.A(\_116_[25] ),
    .B(_05687_),
    .Y(_05688_));
 sky130_fd_sc_hd__o21ai_1 _11662_ (.A1(_05680_),
    .A2(_05683_),
    .B1(_05678_),
    .Y(_05689_));
 sky130_fd_sc_hd__and2_1 _11663_ (.A(_05688_),
    .B(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__o21ai_1 _11664_ (.A1(_05688_),
    .A2(_05689_),
    .B1(_05263_),
    .Y(_05691_));
 sky130_fd_sc_hd__o22a_1 _11665_ (.A1(\_149_[25] ),
    .A2(_05279_),
    .B1(_05690_),
    .B2(_05691_),
    .X(_00780_));
 sky130_fd_sc_hd__xnor2_1 _11666_ (.A(\_118_[29] ),
    .B(\_118_[1] ),
    .Y(_05692_));
 sky130_fd_sc_hd__xnor2_1 _11667_ (.A(\_118_[12] ),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__nand2_1 _11668_ (.A(\_116_[26] ),
    .B(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__or2_1 _11669_ (.A(\_116_[26] ),
    .B(_05693_),
    .X(_05695_));
 sky130_fd_sc_hd__nand2_1 _11670_ (.A(_05694_),
    .B(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__or2_1 _11671_ (.A(_05680_),
    .B(_05688_),
    .X(_05697_));
 sky130_fd_sc_hd__o211a_1 _11672_ (.A1(\_116_[25] ),
    .A2(_05687_),
    .B1(_05677_),
    .C1(\_116_[24] ),
    .X(_05698_));
 sky130_fd_sc_hd__a21oi_1 _11673_ (.A1(\_116_[25] ),
    .A2(_05687_),
    .B1(_05698_),
    .Y(_05699_));
 sky130_fd_sc_hd__o21ai_1 _11674_ (.A1(_05683_),
    .A2(_05697_),
    .B1(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__xnor2_1 _11675_ (.A(_05696_),
    .B(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__mux2_1 _11676_ (.A0(\_149_[26] ),
    .A1(_05701_),
    .S(_05625_),
    .X(_05702_));
 sky130_fd_sc_hd__clkbuf_1 _11677_ (.A(_05702_),
    .X(_00781_));
 sky130_fd_sc_hd__xnor2_1 _11678_ (.A(\_118_[30] ),
    .B(\_118_[2] ),
    .Y(_05703_));
 sky130_fd_sc_hd__xnor2_1 _11679_ (.A(\_118_[13] ),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__nand2_1 _11680_ (.A(\_116_[27] ),
    .B(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hd__or2_1 _11681_ (.A(\_116_[27] ),
    .B(_05704_),
    .X(_05706_));
 sky130_fd_sc_hd__nand2_1 _11682_ (.A(_05705_),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__a21bo_1 _11683_ (.A1(_05695_),
    .A2(_05700_),
    .B1_N(_05694_),
    .X(_05708_));
 sky130_fd_sc_hd__xnor2_1 _11684_ (.A(_05707_),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__mux2_1 _11685_ (.A0(\_149_[27] ),
    .A1(_05709_),
    .S(_05625_),
    .X(_05710_));
 sky130_fd_sc_hd__clkbuf_1 _11686_ (.A(_05710_),
    .X(_00782_));
 sky130_fd_sc_hd__xnor2_1 _11687_ (.A(\_118_[14] ),
    .B(\_118_[31] ),
    .Y(_05711_));
 sky130_fd_sc_hd__xnor2_1 _11688_ (.A(\_118_[3] ),
    .B(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__nand2_1 _11689_ (.A(\_116_[28] ),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__or2_1 _11690_ (.A(\_116_[28] ),
    .B(_05712_),
    .X(_05714_));
 sky130_fd_sc_hd__nand2_1 _11691_ (.A(_05713_),
    .B(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__or2_1 _11692_ (.A(_05696_),
    .B(_05707_),
    .X(_05716_));
 sky130_fd_sc_hd__nor2_1 _11693_ (.A(\_116_[27] ),
    .B(_05704_),
    .Y(_05717_));
 sky130_fd_sc_hd__o221a_1 _11694_ (.A1(_05694_),
    .A2(_05717_),
    .B1(_05716_),
    .B2(_05699_),
    .C1(_05705_),
    .X(_05718_));
 sky130_fd_sc_hd__o31a_1 _11695_ (.A1(_05683_),
    .A2(_05697_),
    .A3(_05716_),
    .B1(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__xor2_1 _11696_ (.A(_05715_),
    .B(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__mux2_1 _11697_ (.A0(\_149_[28] ),
    .A1(_05720_),
    .S(_05625_),
    .X(_05721_));
 sky130_fd_sc_hd__clkbuf_1 _11698_ (.A(_05721_),
    .X(_00783_));
 sky130_fd_sc_hd__or2_1 _11699_ (.A(\_118_[4] ),
    .B(\_118_[15] ),
    .X(_05722_));
 sky130_fd_sc_hd__nand2_1 _11700_ (.A(\_118_[4] ),
    .B(\_118_[15] ),
    .Y(_05723_));
 sky130_fd_sc_hd__a21oi_1 _11701_ (.A1(_05722_),
    .A2(_05723_),
    .B1(\_116_[29] ),
    .Y(_05724_));
 sky130_fd_sc_hd__inv_2 _11702_ (.A(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__nand3_1 _11703_ (.A(\_116_[29] ),
    .B(_05722_),
    .C(_05723_),
    .Y(_05726_));
 sky130_fd_sc_hd__nand2_1 _11704_ (.A(_05725_),
    .B(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__o21ai_1 _11705_ (.A1(_05715_),
    .A2(_05719_),
    .B1(_05713_),
    .Y(_05728_));
 sky130_fd_sc_hd__xnor2_1 _11706_ (.A(_05727_),
    .B(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__mux2_1 _11707_ (.A0(\_149_[29] ),
    .A1(_05729_),
    .S(_05625_),
    .X(_05730_));
 sky130_fd_sc_hd__clkbuf_1 _11708_ (.A(_05730_),
    .X(_00784_));
 sky130_fd_sc_hd__o211ai_2 _11709_ (.A1(_05715_),
    .A2(_05719_),
    .B1(_05726_),
    .C1(_05713_),
    .Y(_05731_));
 sky130_fd_sc_hd__xor2_1 _11710_ (.A(\_118_[5] ),
    .B(\_118_[16] ),
    .X(_05732_));
 sky130_fd_sc_hd__xor2_1 _11711_ (.A(\_116_[30] ),
    .B(_05732_),
    .X(_05733_));
 sky130_fd_sc_hd__and3_1 _11712_ (.A(_05725_),
    .B(_05731_),
    .C(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__a21o_1 _11713_ (.A1(_05725_),
    .A2(_05731_),
    .B1(_05733_),
    .X(_05735_));
 sky130_fd_sc_hd__nand2_1 _11714_ (.A(_05263_),
    .B(_05735_),
    .Y(_05736_));
 sky130_fd_sc_hd__a2bb2o_1 _11715_ (.A1_N(_05734_),
    .A2_N(_05736_),
    .B1(\_149_[30] ),
    .B2(_05262_),
    .X(_00785_));
 sky130_fd_sc_hd__a32o_1 _11716_ (.A1(_05725_),
    .A2(_05731_),
    .A3(_05733_),
    .B1(_05732_),
    .B2(\_116_[30] ),
    .X(_05737_));
 sky130_fd_sc_hd__xor2_1 _11717_ (.A(\_118_[17] ),
    .B(\_116_[31] ),
    .X(_05738_));
 sky130_fd_sc_hd__xnor2_1 _11718_ (.A(\_118_[6] ),
    .B(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__xnor2_1 _11719_ (.A(_05737_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__mux2_1 _11720_ (.A0(\_149_[31] ),
    .A1(_05740_),
    .S(_05625_),
    .X(_05741_));
 sky130_fd_sc_hd__clkbuf_1 _11721_ (.A(_05741_),
    .X(_00786_));
 sky130_fd_sc_hd__buf_4 _11722_ (.A(_01358_),
    .X(_05742_));
 sky130_fd_sc_hd__xnor2_1 _11723_ (.A(\_140_[17] ),
    .B(\_140_[10] ),
    .Y(_05743_));
 sky130_fd_sc_hd__xnor2_1 _11724_ (.A(\_140_[19] ),
    .B(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__nand2_1 _11725_ (.A(\_152_[0] ),
    .B(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__or2_1 _11726_ (.A(\_152_[0] ),
    .B(_05744_),
    .X(_05746_));
 sky130_fd_sc_hd__and2_1 _11727_ (.A(net1),
    .B(_01274_),
    .X(_05747_));
 sky130_fd_sc_hd__a31o_1 _11728_ (.A1(_05742_),
    .A2(_05745_),
    .A3(_05746_),
    .B1(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__mux2_1 _11729_ (.A0(\_142_[0] ),
    .A1(_05748_),
    .S(_05625_),
    .X(_05749_));
 sky130_fd_sc_hd__clkbuf_1 _11730_ (.A(_05749_),
    .X(_00787_));
 sky130_fd_sc_hd__xnor2_1 _11731_ (.A(\_140_[18] ),
    .B(\_140_[11] ),
    .Y(_05750_));
 sky130_fd_sc_hd__xnor2_1 _11732_ (.A(\_140_[20] ),
    .B(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__xnor2_1 _11733_ (.A(\_152_[1] ),
    .B(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__xor2_1 _11734_ (.A(_05745_),
    .B(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__mux2_1 _11735_ (.A0(net12),
    .A1(_05753_),
    .S(_05742_),
    .X(_05754_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(\_142_[1] ),
    .A1(_05754_),
    .S(_05625_),
    .X(_05755_));
 sky130_fd_sc_hd__clkbuf_1 _11737_ (.A(_05755_),
    .X(_00788_));
 sky130_fd_sc_hd__xnor2_1 _11738_ (.A(\_140_[21] ),
    .B(\_140_[12] ),
    .Y(_05756_));
 sky130_fd_sc_hd__xnor2_1 _11739_ (.A(\_140_[19] ),
    .B(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__nand2_1 _11740_ (.A(\_152_[2] ),
    .B(_05757_),
    .Y(_05758_));
 sky130_fd_sc_hd__or2_1 _11741_ (.A(\_152_[2] ),
    .B(_05757_),
    .X(_05759_));
 sky130_fd_sc_hd__nand2_1 _11742_ (.A(_05758_),
    .B(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__nand2_1 _11743_ (.A(\_152_[1] ),
    .B(_05751_),
    .Y(_05761_));
 sky130_fd_sc_hd__o21ai_1 _11744_ (.A1(_05745_),
    .A2(_05752_),
    .B1(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__xnor2_1 _11745_ (.A(_05760_),
    .B(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__mux2_1 _11746_ (.A0(net23),
    .A1(_05763_),
    .S(_05742_),
    .X(_05764_));
 sky130_fd_sc_hd__clkbuf_4 _11747_ (.A(_01361_),
    .X(_05765_));
 sky130_fd_sc_hd__mux2_1 _11748_ (.A0(\_142_[2] ),
    .A1(_05764_),
    .S(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__clkbuf_1 _11749_ (.A(_05766_),
    .X(_00789_));
 sky130_fd_sc_hd__xnor2_1 _11750_ (.A(\_140_[22] ),
    .B(\_140_[13] ),
    .Y(_05767_));
 sky130_fd_sc_hd__xnor2_1 _11751_ (.A(\_140_[20] ),
    .B(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__and2_1 _11752_ (.A(\_152_[3] ),
    .B(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__or2_1 _11753_ (.A(\_152_[3] ),
    .B(_05768_),
    .X(_05770_));
 sky130_fd_sc_hd__or2b_1 _11754_ (.A(_05769_),
    .B_N(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__a21bo_1 _11755_ (.A1(_05759_),
    .A2(_05762_),
    .B1_N(_05758_),
    .X(_05772_));
 sky130_fd_sc_hd__xnor2_1 _11756_ (.A(_05771_),
    .B(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__mux2_1 _11757_ (.A0(net26),
    .A1(_05773_),
    .S(_05742_),
    .X(_05774_));
 sky130_fd_sc_hd__mux2_1 _11758_ (.A0(\_142_[3] ),
    .A1(_05774_),
    .S(_05765_),
    .X(_05775_));
 sky130_fd_sc_hd__clkbuf_1 _11759_ (.A(_05775_),
    .X(_00790_));
 sky130_fd_sc_hd__clkbuf_4 _11760_ (.A(_01274_),
    .X(_05776_));
 sky130_fd_sc_hd__a21o_1 _11761_ (.A1(_05770_),
    .A2(_05772_),
    .B1(_05769_),
    .X(_05777_));
 sky130_fd_sc_hd__xnor2_1 _11762_ (.A(\_140_[23] ),
    .B(\_140_[14] ),
    .Y(_05778_));
 sky130_fd_sc_hd__xnor2_1 _11763_ (.A(\_140_[21] ),
    .B(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__nand2_1 _11764_ (.A(\_152_[4] ),
    .B(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__or2_1 _11765_ (.A(\_152_[4] ),
    .B(_05779_),
    .X(_05781_));
 sky130_fd_sc_hd__nand2_1 _11766_ (.A(_05780_),
    .B(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__inv_2 _11767_ (.A(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__or2_1 _11768_ (.A(_05777_),
    .B(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__clkbuf_4 _11769_ (.A(_01358_),
    .X(_05785_));
 sky130_fd_sc_hd__nand2_1 _11770_ (.A(_05777_),
    .B(_05783_),
    .Y(_05786_));
 sky130_fd_sc_hd__and2_1 _11771_ (.A(_05785_),
    .B(_05786_),
    .X(_05787_));
 sky130_fd_sc_hd__a22o_1 _11772_ (.A1(net27),
    .A2(_05776_),
    .B1(_05784_),
    .B2(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__mux2_1 _11773_ (.A0(\_142_[4] ),
    .A1(_05788_),
    .S(_05765_),
    .X(_05789_));
 sky130_fd_sc_hd__clkbuf_1 _11774_ (.A(_05789_),
    .X(_00791_));
 sky130_fd_sc_hd__xnor2_1 _11775_ (.A(\_140_[24] ),
    .B(\_140_[15] ),
    .Y(_05790_));
 sky130_fd_sc_hd__xnor2_1 _11776_ (.A(\_140_[22] ),
    .B(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__nand2_1 _11777_ (.A(\_152_[5] ),
    .B(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__nor2_1 _11778_ (.A(\_152_[5] ),
    .B(_05791_),
    .Y(_05793_));
 sky130_fd_sc_hd__inv_2 _11779_ (.A(_05793_),
    .Y(_05794_));
 sky130_fd_sc_hd__nand2_1 _11780_ (.A(_05792_),
    .B(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__a21oi_1 _11781_ (.A1(_05780_),
    .A2(_05786_),
    .B1(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__a31o_1 _11782_ (.A1(_05780_),
    .A2(_05786_),
    .A3(_05795_),
    .B1(_01274_),
    .X(_05797_));
 sky130_fd_sc_hd__a2bb2o_1 _11783_ (.A1_N(_05796_),
    .A2_N(_05797_),
    .B1(net28),
    .B2(_05776_),
    .X(_05798_));
 sky130_fd_sc_hd__mux2_1 _11784_ (.A0(\_142_[5] ),
    .A1(_05798_),
    .S(_05765_),
    .X(_05799_));
 sky130_fd_sc_hd__clkbuf_1 _11785_ (.A(_05799_),
    .X(_00792_));
 sky130_fd_sc_hd__nand2_1 _11786_ (.A(_05780_),
    .B(_05792_),
    .Y(_05800_));
 sky130_fd_sc_hd__a21oi_1 _11787_ (.A1(_05777_),
    .A2(_05783_),
    .B1(_05800_),
    .Y(_05801_));
 sky130_fd_sc_hd__xnor2_1 _11788_ (.A(\_140_[25] ),
    .B(\_140_[16] ),
    .Y(_05802_));
 sky130_fd_sc_hd__xnor2_1 _11789_ (.A(\_140_[23] ),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__nand2_1 _11790_ (.A(\_152_[6] ),
    .B(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__or2_1 _11791_ (.A(\_152_[6] ),
    .B(_05803_),
    .X(_05805_));
 sky130_fd_sc_hd__nand2_1 _11792_ (.A(_05804_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__o21ai_1 _11793_ (.A1(_05793_),
    .A2(_05801_),
    .B1(_05806_),
    .Y(_05807_));
 sky130_fd_sc_hd__or3_1 _11794_ (.A(_05793_),
    .B(_05806_),
    .C(_05801_),
    .X(_05808_));
 sky130_fd_sc_hd__and2_1 _11795_ (.A(_01358_),
    .B(_05808_),
    .X(_05809_));
 sky130_fd_sc_hd__a22o_1 _11796_ (.A1(net29),
    .A2(_05776_),
    .B1(_05807_),
    .B2(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__mux2_1 _11797_ (.A0(\_142_[6] ),
    .A1(_05810_),
    .S(_05765_),
    .X(_05811_));
 sky130_fd_sc_hd__clkbuf_1 _11798_ (.A(_05811_),
    .X(_00793_));
 sky130_fd_sc_hd__xnor2_1 _11799_ (.A(\_140_[24] ),
    .B(\_140_[26] ),
    .Y(_05812_));
 sky130_fd_sc_hd__xnor2_1 _11800_ (.A(\_140_[17] ),
    .B(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__nand2_1 _11801_ (.A(\_152_[7] ),
    .B(_05813_),
    .Y(_05814_));
 sky130_fd_sc_hd__nor2_1 _11802_ (.A(\_152_[7] ),
    .B(_05813_),
    .Y(_05815_));
 sky130_fd_sc_hd__inv_2 _11803_ (.A(_05815_),
    .Y(_05816_));
 sky130_fd_sc_hd__nand2_1 _11804_ (.A(_05814_),
    .B(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__a21o_1 _11805_ (.A1(_05804_),
    .A2(_05808_),
    .B1(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__a31oi_1 _11806_ (.A1(_05804_),
    .A2(_05808_),
    .A3(_05817_),
    .B1(_05776_),
    .Y(_05819_));
 sky130_fd_sc_hd__a221o_1 _11807_ (.A1(net30),
    .A2(_05776_),
    .B1(_05818_),
    .B2(_05819_),
    .C1(_01368_),
    .X(_05820_));
 sky130_fd_sc_hd__o21a_1 _11808_ (.A1(\_142_[7] ),
    .A2(_05279_),
    .B1(_05820_),
    .X(_00794_));
 sky130_fd_sc_hd__xnor2_1 _11809_ (.A(\_140_[25] ),
    .B(\_140_[27] ),
    .Y(_05821_));
 sky130_fd_sc_hd__xnor2_1 _11810_ (.A(\_140_[18] ),
    .B(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__nand2_1 _11811_ (.A(\_152_[8] ),
    .B(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__or2_1 _11812_ (.A(\_152_[8] ),
    .B(_05822_),
    .X(_05824_));
 sky130_fd_sc_hd__nand2_1 _11813_ (.A(_05823_),
    .B(_05824_),
    .Y(_05825_));
 sky130_fd_sc_hd__and2_1 _11814_ (.A(_05804_),
    .B(_05814_),
    .X(_05826_));
 sky130_fd_sc_hd__o31a_1 _11815_ (.A1(_05793_),
    .A2(_05806_),
    .A3(_05801_),
    .B1(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__or2_1 _11816_ (.A(_05815_),
    .B(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__nand2_1 _11817_ (.A(_05825_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__or2_1 _11818_ (.A(_05825_),
    .B(_05828_),
    .X(_05830_));
 sky130_fd_sc_hd__and3_1 _11819_ (.A(_05742_),
    .B(_05829_),
    .C(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__a211o_1 _11820_ (.A1(net31),
    .A2(_05776_),
    .B1(_01368_),
    .C1(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__o21a_1 _11821_ (.A1(\_142_[8] ),
    .A2(_05279_),
    .B1(_05832_),
    .X(_00795_));
 sky130_fd_sc_hd__xnor2_1 _11822_ (.A(\_140_[26] ),
    .B(\_140_[28] ),
    .Y(_05833_));
 sky130_fd_sc_hd__xnor2_1 _11823_ (.A(\_140_[19] ),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__nand2_1 _11824_ (.A(\_152_[9] ),
    .B(_05834_),
    .Y(_05835_));
 sky130_fd_sc_hd__nor2_1 _11825_ (.A(\_152_[9] ),
    .B(_05834_),
    .Y(_05836_));
 sky130_fd_sc_hd__inv_2 _11826_ (.A(_05836_),
    .Y(_05837_));
 sky130_fd_sc_hd__nand2_1 _11827_ (.A(_05835_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__a21oi_1 _11828_ (.A1(_05823_),
    .A2(_05830_),
    .B1(_05838_),
    .Y(_05839_));
 sky130_fd_sc_hd__a31o_1 _11829_ (.A1(_05823_),
    .A2(_05830_),
    .A3(_05838_),
    .B1(_01274_),
    .X(_05840_));
 sky130_fd_sc_hd__a2bb2o_1 _11830_ (.A1_N(_05839_),
    .A2_N(_05840_),
    .B1(net32),
    .B2(_05776_),
    .X(_05841_));
 sky130_fd_sc_hd__mux2_1 _11831_ (.A0(\_142_[9] ),
    .A1(_05841_),
    .S(_05765_),
    .X(_05842_));
 sky130_fd_sc_hd__clkbuf_1 _11832_ (.A(_05842_),
    .X(_00796_));
 sky130_fd_sc_hd__xnor2_1 _11833_ (.A(\_140_[27] ),
    .B(\_140_[29] ),
    .Y(_05843_));
 sky130_fd_sc_hd__xnor2_1 _11834_ (.A(\_140_[20] ),
    .B(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__nand2_1 _11835_ (.A(\_152_[10] ),
    .B(_05844_),
    .Y(_05845_));
 sky130_fd_sc_hd__or2_1 _11836_ (.A(\_152_[10] ),
    .B(_05844_),
    .X(_05846_));
 sky130_fd_sc_hd__nand2_1 _11837_ (.A(_05845_),
    .B(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__and2_1 _11838_ (.A(_05823_),
    .B(_05835_),
    .X(_05848_));
 sky130_fd_sc_hd__o31a_1 _11839_ (.A1(_05815_),
    .A2(_05825_),
    .A3(_05827_),
    .B1(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__or2_1 _11840_ (.A(_05836_),
    .B(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__xor2_1 _11841_ (.A(_05847_),
    .B(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__buf_4 _11842_ (.A(_01358_),
    .X(_05852_));
 sky130_fd_sc_hd__mux2_1 _11843_ (.A0(net2),
    .A1(_05851_),
    .S(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__mux2_1 _11844_ (.A0(\_142_[10] ),
    .A1(_05853_),
    .S(_05765_),
    .X(_05854_));
 sky130_fd_sc_hd__clkbuf_1 _11845_ (.A(_05854_),
    .X(_00797_));
 sky130_fd_sc_hd__xnor2_1 _11846_ (.A(\_140_[28] ),
    .B(\_140_[30] ),
    .Y(_05855_));
 sky130_fd_sc_hd__xnor2_1 _11847_ (.A(\_140_[21] ),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__and2_1 _11848_ (.A(\_152_[11] ),
    .B(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__or2_1 _11849_ (.A(\_152_[11] ),
    .B(_05856_),
    .X(_05858_));
 sky130_fd_sc_hd__or2b_1 _11850_ (.A(_05857_),
    .B_N(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__o31ai_2 _11851_ (.A1(_05836_),
    .A2(_05847_),
    .A3(_05849_),
    .B1(_05845_),
    .Y(_05860_));
 sky130_fd_sc_hd__xnor2_1 _11852_ (.A(_05859_),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__mux2_1 _11853_ (.A0(net3),
    .A1(_05861_),
    .S(_05852_),
    .X(_05862_));
 sky130_fd_sc_hd__mux2_1 _11854_ (.A0(\_142_[11] ),
    .A1(_05862_),
    .S(_05765_),
    .X(_05863_));
 sky130_fd_sc_hd__clkbuf_1 _11855_ (.A(_05863_),
    .X(_00798_));
 sky130_fd_sc_hd__a21oi_2 _11856_ (.A1(_05858_),
    .A2(_05860_),
    .B1(_05857_),
    .Y(_05864_));
 sky130_fd_sc_hd__xnor2_1 _11857_ (.A(\_140_[29] ),
    .B(\_140_[31] ),
    .Y(_05865_));
 sky130_fd_sc_hd__xnor2_1 _11858_ (.A(\_140_[22] ),
    .B(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__nand2_1 _11859_ (.A(\_152_[12] ),
    .B(_05866_),
    .Y(_05867_));
 sky130_fd_sc_hd__or2_1 _11860_ (.A(\_152_[12] ),
    .B(_05866_),
    .X(_05868_));
 sky130_fd_sc_hd__nand2_1 _11861_ (.A(_05867_),
    .B(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__nand2_1 _11862_ (.A(_05864_),
    .B(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__o21a_1 _11863_ (.A1(_05864_),
    .A2(_05869_),
    .B1(_05785_),
    .X(_05871_));
 sky130_fd_sc_hd__a22o_1 _11864_ (.A1(net4),
    .A2(_05776_),
    .B1(_05870_),
    .B2(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(\_142_[12] ),
    .A1(_05872_),
    .S(_05765_),
    .X(_05873_));
 sky130_fd_sc_hd__clkbuf_1 _11866_ (.A(_05873_),
    .X(_00799_));
 sky130_fd_sc_hd__xnor2_1 _11867_ (.A(\_140_[30] ),
    .B(\_140_[0] ),
    .Y(_05874_));
 sky130_fd_sc_hd__xnor2_1 _11868_ (.A(\_140_[23] ),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__nand2_1 _11869_ (.A(\_152_[13] ),
    .B(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__nor2_1 _11870_ (.A(\_152_[13] ),
    .B(_05875_),
    .Y(_05877_));
 sky130_fd_sc_hd__inv_2 _11871_ (.A(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__nand2_1 _11872_ (.A(_05876_),
    .B(_05878_),
    .Y(_05879_));
 sky130_fd_sc_hd__o21ai_1 _11873_ (.A1(_05864_),
    .A2(_05869_),
    .B1(_05867_),
    .Y(_05880_));
 sky130_fd_sc_hd__xnor2_1 _11874_ (.A(_05879_),
    .B(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__mux2_1 _11875_ (.A0(net5),
    .A1(_05881_),
    .S(_05852_),
    .X(_05882_));
 sky130_fd_sc_hd__mux2_1 _11876_ (.A0(\_142_[13] ),
    .A1(_05882_),
    .S(_05765_),
    .X(_05883_));
 sky130_fd_sc_hd__clkbuf_1 _11877_ (.A(_05883_),
    .X(_00800_));
 sky130_fd_sc_hd__xnor2_2 _11878_ (.A(\_140_[31] ),
    .B(\_140_[1] ),
    .Y(_05884_));
 sky130_fd_sc_hd__xnor2_2 _11879_ (.A(\_140_[24] ),
    .B(_05884_),
    .Y(_05885_));
 sky130_fd_sc_hd__nand2_1 _11880_ (.A(\_152_[14] ),
    .B(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__or2_1 _11881_ (.A(\_152_[14] ),
    .B(_05885_),
    .X(_05887_));
 sky130_fd_sc_hd__nand2_1 _11882_ (.A(_05886_),
    .B(_05887_),
    .Y(_05888_));
 sky130_fd_sc_hd__a21o_1 _11883_ (.A1(_05867_),
    .A2(_05876_),
    .B1(_05877_),
    .X(_05889_));
 sky130_fd_sc_hd__o31a_2 _11884_ (.A1(_05864_),
    .A2(_05869_),
    .A3(_05879_),
    .B1(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__xor2_1 _11885_ (.A(_05888_),
    .B(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__mux2_1 _11886_ (.A0(net6),
    .A1(_05891_),
    .S(_05852_),
    .X(_05892_));
 sky130_fd_sc_hd__clkbuf_4 _11887_ (.A(_01361_),
    .X(_05893_));
 sky130_fd_sc_hd__mux2_1 _11888_ (.A0(\_142_[14] ),
    .A1(_05892_),
    .S(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__clkbuf_1 _11889_ (.A(_05894_),
    .X(_00801_));
 sky130_fd_sc_hd__xnor2_2 _11890_ (.A(\_140_[0] ),
    .B(\_140_[2] ),
    .Y(_05895_));
 sky130_fd_sc_hd__xnor2_2 _11891_ (.A(\_140_[25] ),
    .B(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__xnor2_1 _11892_ (.A(\_152_[15] ),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__o21ai_1 _11893_ (.A1(_05888_),
    .A2(_05890_),
    .B1(_05886_),
    .Y(_05898_));
 sky130_fd_sc_hd__xnor2_1 _11894_ (.A(_05897_),
    .B(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__mux2_1 _11895_ (.A0(net7),
    .A1(_05899_),
    .S(_05852_),
    .X(_05900_));
 sky130_fd_sc_hd__mux2_1 _11896_ (.A0(\_142_[15] ),
    .A1(_05900_),
    .S(_05893_),
    .X(_05901_));
 sky130_fd_sc_hd__clkbuf_1 _11897_ (.A(_05901_),
    .X(_00802_));
 sky130_fd_sc_hd__xnor2_2 _11898_ (.A(\_140_[1] ),
    .B(\_140_[3] ),
    .Y(_05902_));
 sky130_fd_sc_hd__xnor2_2 _11899_ (.A(\_140_[26] ),
    .B(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__nand2_1 _11900_ (.A(\_152_[16] ),
    .B(_05903_),
    .Y(_05904_));
 sky130_fd_sc_hd__or2_1 _11901_ (.A(\_152_[16] ),
    .B(_05903_),
    .X(_05905_));
 sky130_fd_sc_hd__nand2_1 _11902_ (.A(_05904_),
    .B(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__a22o_1 _11903_ (.A1(\_152_[14] ),
    .A2(_05885_),
    .B1(_05896_),
    .B2(\_152_[15] ),
    .X(_05907_));
 sky130_fd_sc_hd__o21ai_1 _11904_ (.A1(\_152_[15] ),
    .A2(_05896_),
    .B1(_05907_),
    .Y(_05908_));
 sky130_fd_sc_hd__o31a_2 _11905_ (.A1(_05888_),
    .A2(_05890_),
    .A3(_05897_),
    .B1(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__xor2_1 _11906_ (.A(_05906_),
    .B(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__mux2_1 _11907_ (.A0(net8),
    .A1(_05910_),
    .S(_05852_),
    .X(_05911_));
 sky130_fd_sc_hd__mux2_1 _11908_ (.A0(\_142_[16] ),
    .A1(_05911_),
    .S(_05893_),
    .X(_05912_));
 sky130_fd_sc_hd__clkbuf_1 _11909_ (.A(_05912_),
    .X(_00803_));
 sky130_fd_sc_hd__xnor2_2 _11910_ (.A(\_140_[2] ),
    .B(\_140_[4] ),
    .Y(_05913_));
 sky130_fd_sc_hd__xnor2_2 _11911_ (.A(\_140_[27] ),
    .B(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__xnor2_1 _11912_ (.A(\_152_[17] ),
    .B(_05914_),
    .Y(_05915_));
 sky130_fd_sc_hd__o21ai_1 _11913_ (.A1(_05906_),
    .A2(_05909_),
    .B1(_05904_),
    .Y(_05916_));
 sky130_fd_sc_hd__xnor2_1 _11914_ (.A(_05915_),
    .B(_05916_),
    .Y(_05917_));
 sky130_fd_sc_hd__mux2_1 _11915_ (.A0(net9),
    .A1(_05917_),
    .S(_05852_),
    .X(_05918_));
 sky130_fd_sc_hd__mux2_1 _11916_ (.A0(\_142_[17] ),
    .A1(_05918_),
    .S(_05893_),
    .X(_05919_));
 sky130_fd_sc_hd__clkbuf_1 _11917_ (.A(_05919_),
    .X(_00804_));
 sky130_fd_sc_hd__xnor2_1 _11918_ (.A(\_140_[3] ),
    .B(\_140_[5] ),
    .Y(_05920_));
 sky130_fd_sc_hd__xnor2_1 _11919_ (.A(\_140_[28] ),
    .B(_05920_),
    .Y(_05921_));
 sky130_fd_sc_hd__nand2_1 _11920_ (.A(\_152_[18] ),
    .B(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__or2_1 _11921_ (.A(\_152_[18] ),
    .B(_05921_),
    .X(_05923_));
 sky130_fd_sc_hd__nand2_1 _11922_ (.A(_05922_),
    .B(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__or2_1 _11923_ (.A(_05906_),
    .B(_05915_),
    .X(_05925_));
 sky130_fd_sc_hd__o211a_1 _11924_ (.A1(\_152_[17] ),
    .A2(_05914_),
    .B1(_05903_),
    .C1(\_152_[16] ),
    .X(_05926_));
 sky130_fd_sc_hd__a21oi_1 _11925_ (.A1(\_152_[17] ),
    .A2(_05914_),
    .B1(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__o21a_1 _11926_ (.A1(_05909_),
    .A2(_05925_),
    .B1(_05927_),
    .X(_05928_));
 sky130_fd_sc_hd__xor2_1 _11927_ (.A(_05924_),
    .B(_05928_),
    .X(_05929_));
 sky130_fd_sc_hd__mux2_1 _11928_ (.A0(net10),
    .A1(_05929_),
    .S(_05852_),
    .X(_05930_));
 sky130_fd_sc_hd__mux2_1 _11929_ (.A0(\_142_[18] ),
    .A1(_05930_),
    .S(_05893_),
    .X(_05931_));
 sky130_fd_sc_hd__clkbuf_1 _11930_ (.A(_05931_),
    .X(_00805_));
 sky130_fd_sc_hd__xnor2_2 _11931_ (.A(\_140_[4] ),
    .B(\_140_[6] ),
    .Y(_05932_));
 sky130_fd_sc_hd__xnor2_2 _11932_ (.A(\_140_[29] ),
    .B(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__nand2_1 _11933_ (.A(\_152_[19] ),
    .B(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__or2_1 _11934_ (.A(\_152_[19] ),
    .B(_05933_),
    .X(_05935_));
 sky130_fd_sc_hd__nand2_1 _11935_ (.A(_05934_),
    .B(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__o21ai_1 _11936_ (.A1(_05924_),
    .A2(_05928_),
    .B1(_05922_),
    .Y(_05937_));
 sky130_fd_sc_hd__and2_1 _11937_ (.A(_05936_),
    .B(_05937_),
    .X(_05938_));
 sky130_fd_sc_hd__o21ai_1 _11938_ (.A1(_05936_),
    .A2(_05937_),
    .B1(_05785_),
    .Y(_05939_));
 sky130_fd_sc_hd__o22a_1 _11939_ (.A1(net11),
    .A2(_05742_),
    .B1(_05938_),
    .B2(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__mux2_1 _11940_ (.A0(\_142_[19] ),
    .A1(_05940_),
    .S(_05893_),
    .X(_05941_));
 sky130_fd_sc_hd__clkbuf_1 _11941_ (.A(_05941_),
    .X(_00806_));
 sky130_fd_sc_hd__xnor2_1 _11942_ (.A(\_140_[5] ),
    .B(\_140_[7] ),
    .Y(_05942_));
 sky130_fd_sc_hd__xnor2_1 _11943_ (.A(\_140_[30] ),
    .B(_05942_),
    .Y(_05943_));
 sky130_fd_sc_hd__nand2_1 _11944_ (.A(\_152_[20] ),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__or2_1 _11945_ (.A(\_152_[20] ),
    .B(_05943_),
    .X(_05945_));
 sky130_fd_sc_hd__nand2_1 _11946_ (.A(_05944_),
    .B(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__or2_1 _11947_ (.A(_05924_),
    .B(_05936_),
    .X(_05947_));
 sky130_fd_sc_hd__or2_1 _11948_ (.A(_05925_),
    .B(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__nor2_1 _11949_ (.A(\_152_[19] ),
    .B(_05933_),
    .Y(_05949_));
 sky130_fd_sc_hd__o221a_1 _11950_ (.A1(_05922_),
    .A2(_05949_),
    .B1(_05947_),
    .B2(_05927_),
    .C1(_05934_),
    .X(_05950_));
 sky130_fd_sc_hd__o21a_1 _11951_ (.A1(_05909_),
    .A2(_05948_),
    .B1(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__xor2_1 _11952_ (.A(_05946_),
    .B(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__mux2_1 _11953_ (.A0(net13),
    .A1(_05952_),
    .S(_05852_),
    .X(_05953_));
 sky130_fd_sc_hd__mux2_1 _11954_ (.A0(\_142_[20] ),
    .A1(_05953_),
    .S(_05893_),
    .X(_05954_));
 sky130_fd_sc_hd__clkbuf_1 _11955_ (.A(_05954_),
    .X(_00807_));
 sky130_fd_sc_hd__or2_1 _11956_ (.A(_05946_),
    .B(_05951_),
    .X(_05955_));
 sky130_fd_sc_hd__nand2_1 _11957_ (.A(_05944_),
    .B(_05955_),
    .Y(_05956_));
 sky130_fd_sc_hd__xnor2_1 _11958_ (.A(\_140_[6] ),
    .B(\_140_[8] ),
    .Y(_05957_));
 sky130_fd_sc_hd__xnor2_2 _11959_ (.A(\_140_[31] ),
    .B(_05957_),
    .Y(_05958_));
 sky130_fd_sc_hd__nor2_1 _11960_ (.A(\_152_[21] ),
    .B(_05958_),
    .Y(_05959_));
 sky130_fd_sc_hd__nand2_1 _11961_ (.A(\_152_[21] ),
    .B(_05958_),
    .Y(_05960_));
 sky130_fd_sc_hd__or2b_1 _11962_ (.A(_05959_),
    .B_N(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__xnor2_1 _11963_ (.A(_05956_),
    .B(_05961_),
    .Y(_05962_));
 sky130_fd_sc_hd__mux2_1 _11964_ (.A0(net14),
    .A1(_05962_),
    .S(_05852_),
    .X(_05963_));
 sky130_fd_sc_hd__mux2_1 _11965_ (.A0(\_142_[21] ),
    .A1(_05963_),
    .S(_05893_),
    .X(_05964_));
 sky130_fd_sc_hd__clkbuf_1 _11966_ (.A(_05964_),
    .X(_00808_));
 sky130_fd_sc_hd__xor2_2 _11967_ (.A(\_140_[7] ),
    .B(\_140_[9] ),
    .X(_05965_));
 sky130_fd_sc_hd__nand2_1 _11968_ (.A(\_152_[22] ),
    .B(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__or2_1 _11969_ (.A(\_152_[22] ),
    .B(_05965_),
    .X(_05967_));
 sky130_fd_sc_hd__nand2_1 _11970_ (.A(_05966_),
    .B(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__a21oi_1 _11971_ (.A1(_05944_),
    .A2(_05960_),
    .B1(_05959_),
    .Y(_05969_));
 sky130_fd_sc_hd__o21bai_1 _11972_ (.A1(_05955_),
    .A2(_05961_),
    .B1_N(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__xnor2_1 _11973_ (.A(_05968_),
    .B(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__or2_1 _11974_ (.A(net15),
    .B(_05742_),
    .X(_05972_));
 sky130_fd_sc_hd__o211a_1 _11975_ (.A1(_05776_),
    .A2(_05971_),
    .B1(_05972_),
    .C1(_05263_),
    .X(_05973_));
 sky130_fd_sc_hd__a21o_1 _11976_ (.A1(\_142_[22] ),
    .A2(_05262_),
    .B1(_05973_),
    .X(_00809_));
 sky130_fd_sc_hd__or2_1 _11977_ (.A(\_140_[10] ),
    .B(\_140_[8] ),
    .X(_05974_));
 sky130_fd_sc_hd__nand2_1 _11978_ (.A(\_140_[10] ),
    .B(\_140_[8] ),
    .Y(_05975_));
 sky130_fd_sc_hd__a21oi_1 _11979_ (.A1(_05974_),
    .A2(_05975_),
    .B1(\_152_[23] ),
    .Y(_05976_));
 sky130_fd_sc_hd__nand3_1 _11980_ (.A(\_152_[23] ),
    .B(_05974_),
    .C(_05975_),
    .Y(_05977_));
 sky130_fd_sc_hd__or2b_1 _11981_ (.A(_05976_),
    .B_N(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__a21bo_1 _11982_ (.A1(_05967_),
    .A2(_05970_),
    .B1_N(_05966_),
    .X(_05979_));
 sky130_fd_sc_hd__xnor2_1 _11983_ (.A(_05978_),
    .B(_05979_),
    .Y(_05980_));
 sky130_fd_sc_hd__mux2_1 _11984_ (.A0(net16),
    .A1(_05980_),
    .S(_05785_),
    .X(_05981_));
 sky130_fd_sc_hd__mux2_1 _11985_ (.A0(\_142_[23] ),
    .A1(_05981_),
    .S(_05893_),
    .X(_05982_));
 sky130_fd_sc_hd__clkbuf_1 _11986_ (.A(_05982_),
    .X(_00810_));
 sky130_fd_sc_hd__xor2_1 _11987_ (.A(\_140_[11] ),
    .B(\_140_[9] ),
    .X(_05983_));
 sky130_fd_sc_hd__nand2_1 _11988_ (.A(\_152_[24] ),
    .B(_05983_),
    .Y(_05984_));
 sky130_fd_sc_hd__or2_1 _11989_ (.A(\_152_[24] ),
    .B(_05983_),
    .X(_05985_));
 sky130_fd_sc_hd__nand2_1 _11990_ (.A(_05984_),
    .B(_05985_),
    .Y(_05986_));
 sky130_fd_sc_hd__nor2_1 _11991_ (.A(_05968_),
    .B(_05978_),
    .Y(_05987_));
 sky130_fd_sc_hd__or3b_1 _11992_ (.A(_05946_),
    .B(_05961_),
    .C_N(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__o2bb2a_1 _11993_ (.A1_N(_05969_),
    .A2_N(_05987_),
    .B1(_05988_),
    .B2(_05950_),
    .X(_05989_));
 sky130_fd_sc_hd__o211a_1 _11994_ (.A1(_05966_),
    .A2(_05976_),
    .B1(_05977_),
    .C1(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__o31a_1 _11995_ (.A1(_05909_),
    .A2(_05948_),
    .A3(_05988_),
    .B1(_05990_),
    .X(_05991_));
 sky130_fd_sc_hd__xor2_1 _11996_ (.A(_05986_),
    .B(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__mux2_1 _11997_ (.A0(net17),
    .A1(_05992_),
    .S(_05785_),
    .X(_05993_));
 sky130_fd_sc_hd__mux2_1 _11998_ (.A0(\_142_[24] ),
    .A1(_05993_),
    .S(_05893_),
    .X(_05994_));
 sky130_fd_sc_hd__clkbuf_1 _11999_ (.A(_05994_),
    .X(_00811_));
 sky130_fd_sc_hd__or2_1 _12000_ (.A(\_140_[10] ),
    .B(\_140_[12] ),
    .X(_05995_));
 sky130_fd_sc_hd__nand2_1 _12001_ (.A(\_140_[10] ),
    .B(\_140_[12] ),
    .Y(_05996_));
 sky130_fd_sc_hd__and3_1 _12002_ (.A(\_152_[25] ),
    .B(_05995_),
    .C(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__a21oi_1 _12003_ (.A1(_05995_),
    .A2(_05996_),
    .B1(\_152_[25] ),
    .Y(_05998_));
 sky130_fd_sc_hd__or2_1 _12004_ (.A(_05997_),
    .B(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__o21ai_1 _12005_ (.A1(_05986_),
    .A2(_05991_),
    .B1(_05984_),
    .Y(_06000_));
 sky130_fd_sc_hd__and2_1 _12006_ (.A(_05999_),
    .B(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__o21ai_1 _12007_ (.A1(_05999_),
    .A2(_06000_),
    .B1(_05785_),
    .Y(_06002_));
 sky130_fd_sc_hd__o22a_1 _12008_ (.A1(net18),
    .A2(_05742_),
    .B1(_06001_),
    .B2(_06002_),
    .X(_06003_));
 sky130_fd_sc_hd__buf_6 _12009_ (.A(_01360_),
    .X(_06004_));
 sky130_fd_sc_hd__buf_4 _12010_ (.A(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__mux2_1 _12011_ (.A0(\_142_[25] ),
    .A1(_06003_),
    .S(_06005_),
    .X(_06006_));
 sky130_fd_sc_hd__clkbuf_1 _12012_ (.A(_06006_),
    .X(_00812_));
 sky130_fd_sc_hd__xor2_1 _12013_ (.A(\_140_[11] ),
    .B(\_140_[13] ),
    .X(_06007_));
 sky130_fd_sc_hd__nand2_1 _12014_ (.A(\_152_[26] ),
    .B(_06007_),
    .Y(_06008_));
 sky130_fd_sc_hd__or2_1 _12015_ (.A(\_152_[26] ),
    .B(_06007_),
    .X(_06009_));
 sky130_fd_sc_hd__nand2_1 _12016_ (.A(_06008_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__or2_1 _12017_ (.A(_05986_),
    .B(_05999_),
    .X(_06011_));
 sky130_fd_sc_hd__nand3_1 _12018_ (.A(\_152_[25] ),
    .B(_05995_),
    .C(_05996_),
    .Y(_06012_));
 sky130_fd_sc_hd__o21a_1 _12019_ (.A1(_05984_),
    .A2(_05998_),
    .B1(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__o21a_1 _12020_ (.A1(_05991_),
    .A2(_06011_),
    .B1(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__xor2_1 _12021_ (.A(_06010_),
    .B(_06014_),
    .X(_06015_));
 sky130_fd_sc_hd__mux2_1 _12022_ (.A0(net19),
    .A1(_06015_),
    .S(_05785_),
    .X(_06016_));
 sky130_fd_sc_hd__mux2_1 _12023_ (.A0(\_142_[26] ),
    .A1(_06016_),
    .S(_06005_),
    .X(_06017_));
 sky130_fd_sc_hd__clkbuf_1 _12024_ (.A(_06017_),
    .X(_00813_));
 sky130_fd_sc_hd__or2_1 _12025_ (.A(\_140_[12] ),
    .B(\_140_[14] ),
    .X(_06018_));
 sky130_fd_sc_hd__nand2_1 _12026_ (.A(\_140_[12] ),
    .B(\_140_[14] ),
    .Y(_06019_));
 sky130_fd_sc_hd__and3_1 _12027_ (.A(\_152_[27] ),
    .B(_06018_),
    .C(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__a21oi_1 _12028_ (.A1(_06018_),
    .A2(_06019_),
    .B1(\_152_[27] ),
    .Y(_06021_));
 sky130_fd_sc_hd__or2_1 _12029_ (.A(_06020_),
    .B(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__o21ai_1 _12030_ (.A1(_06010_),
    .A2(_06014_),
    .B1(_06008_),
    .Y(_06023_));
 sky130_fd_sc_hd__xnor2_1 _12031_ (.A(_06022_),
    .B(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__mux2_1 _12032_ (.A0(net20),
    .A1(_06024_),
    .S(_05785_),
    .X(_06025_));
 sky130_fd_sc_hd__mux2_1 _12033_ (.A0(\_142_[27] ),
    .A1(_06025_),
    .S(_06005_),
    .X(_06026_));
 sky130_fd_sc_hd__clkbuf_1 _12034_ (.A(_06026_),
    .X(_00814_));
 sky130_fd_sc_hd__or3_1 _12035_ (.A(_06010_),
    .B(_06011_),
    .C(_06022_),
    .X(_06027_));
 sky130_fd_sc_hd__o21ba_1 _12036_ (.A1(_06008_),
    .A2(_06021_),
    .B1_N(_06020_),
    .X(_06028_));
 sky130_fd_sc_hd__o31a_1 _12037_ (.A1(_06010_),
    .A2(_06013_),
    .A3(_06022_),
    .B1(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__o21ai_1 _12038_ (.A1(_05991_),
    .A2(_06027_),
    .B1(_06029_),
    .Y(_06030_));
 sky130_fd_sc_hd__xor2_1 _12039_ (.A(\_140_[13] ),
    .B(\_140_[15] ),
    .X(_06031_));
 sky130_fd_sc_hd__and2_1 _12040_ (.A(\_152_[28] ),
    .B(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__nor2_1 _12041_ (.A(\_152_[28] ),
    .B(_06031_),
    .Y(_06033_));
 sky130_fd_sc_hd__nor2_1 _12042_ (.A(_06032_),
    .B(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__xor2_1 _12043_ (.A(_06030_),
    .B(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__mux2_1 _12044_ (.A0(net21),
    .A1(_06035_),
    .S(_05785_),
    .X(_06036_));
 sky130_fd_sc_hd__mux2_1 _12045_ (.A0(\_142_[28] ),
    .A1(_06036_),
    .S(_06005_),
    .X(_06037_));
 sky130_fd_sc_hd__clkbuf_1 _12046_ (.A(_06037_),
    .X(_00815_));
 sky130_fd_sc_hd__a21oi_1 _12047_ (.A1(_06030_),
    .A2(_06034_),
    .B1(_06032_),
    .Y(_06038_));
 sky130_fd_sc_hd__or2_1 _12048_ (.A(\_140_[14] ),
    .B(\_140_[16] ),
    .X(_06039_));
 sky130_fd_sc_hd__nand2_1 _12049_ (.A(\_140_[14] ),
    .B(\_140_[16] ),
    .Y(_06040_));
 sky130_fd_sc_hd__and3_1 _12050_ (.A(\_152_[29] ),
    .B(_06039_),
    .C(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__a21oi_1 _12051_ (.A1(_06039_),
    .A2(_06040_),
    .B1(\_152_[29] ),
    .Y(_06042_));
 sky130_fd_sc_hd__nor2_1 _12052_ (.A(_06041_),
    .B(_06042_),
    .Y(_06043_));
 sky130_fd_sc_hd__xnor2_1 _12053_ (.A(_06038_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__mux2_1 _12054_ (.A0(net22),
    .A1(_06044_),
    .S(_05785_),
    .X(_06045_));
 sky130_fd_sc_hd__mux2_1 _12055_ (.A0(\_142_[29] ),
    .A1(_06045_),
    .S(_06005_),
    .X(_06046_));
 sky130_fd_sc_hd__clkbuf_1 _12056_ (.A(_06046_),
    .X(_00816_));
 sky130_fd_sc_hd__or2_1 _12057_ (.A(\_140_[17] ),
    .B(\_140_[15] ),
    .X(_06047_));
 sky130_fd_sc_hd__nand2_1 _12058_ (.A(\_140_[17] ),
    .B(\_140_[15] ),
    .Y(_06048_));
 sky130_fd_sc_hd__nand3_1 _12059_ (.A(\_152_[30] ),
    .B(_06047_),
    .C(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__a21o_1 _12060_ (.A1(_06047_),
    .A2(_06048_),
    .B1(\_152_[30] ),
    .X(_06050_));
 sky130_fd_sc_hd__nand2_1 _12061_ (.A(_06049_),
    .B(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__inv_2 _12062_ (.A(_06041_),
    .Y(_06052_));
 sky130_fd_sc_hd__a21o_1 _12063_ (.A1(_06038_),
    .A2(_06052_),
    .B1(_06042_),
    .X(_06053_));
 sky130_fd_sc_hd__nand2_1 _12064_ (.A(_06051_),
    .B(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__a211o_1 _12065_ (.A1(_06038_),
    .A2(_06052_),
    .B1(_06042_),
    .C1(_06051_),
    .X(_06055_));
 sky130_fd_sc_hd__and2_1 _12066_ (.A(net24),
    .B(_01274_),
    .X(_06056_));
 sky130_fd_sc_hd__a31o_1 _12067_ (.A1(_05742_),
    .A2(_06054_),
    .A3(_06055_),
    .B1(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__mux2_1 _12068_ (.A0(\_142_[30] ),
    .A1(_06057_),
    .S(_06005_),
    .X(_06058_));
 sky130_fd_sc_hd__clkbuf_1 _12069_ (.A(_06058_),
    .X(_00817_));
 sky130_fd_sc_hd__xnor2_1 _12070_ (.A(\_140_[16] ),
    .B(\_152_[31] ),
    .Y(_06059_));
 sky130_fd_sc_hd__xnor2_1 _12071_ (.A(\_140_[18] ),
    .B(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__a21oi_1 _12072_ (.A1(_06049_),
    .A2(_06055_),
    .B1(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__a311o_1 _12073_ (.A1(_06049_),
    .A2(_06055_),
    .A3(_06060_),
    .B1(_06061_),
    .C1(_05776_),
    .X(_06062_));
 sky130_fd_sc_hd__o21a_1 _12074_ (.A1(net25),
    .A2(_05742_),
    .B1(_05263_),
    .X(_06063_));
 sky130_fd_sc_hd__a22o_1 _12075_ (.A1(\_142_[31] ),
    .A2(_05352_),
    .B1(_06062_),
    .B2(_06063_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _12076_ (.A0(\_140_[0] ),
    .A1(\_142_[0] ),
    .S(_06005_),
    .X(_06064_));
 sky130_fd_sc_hd__clkbuf_1 _12077_ (.A(_06064_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _12078_ (.A0(\_140_[1] ),
    .A1(\_142_[1] ),
    .S(_06005_),
    .X(_06065_));
 sky130_fd_sc_hd__clkbuf_1 _12079_ (.A(_06065_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _12080_ (.A0(\_140_[2] ),
    .A1(\_142_[2] ),
    .S(_06005_),
    .X(_06066_));
 sky130_fd_sc_hd__clkbuf_1 _12081_ (.A(_06066_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _12082_ (.A0(\_140_[3] ),
    .A1(\_142_[3] ),
    .S(_06005_),
    .X(_06067_));
 sky130_fd_sc_hd__clkbuf_1 _12083_ (.A(_06067_),
    .X(_00822_));
 sky130_fd_sc_hd__clkbuf_4 _12084_ (.A(_06004_),
    .X(_06068_));
 sky130_fd_sc_hd__mux2_1 _12085_ (.A0(\_140_[4] ),
    .A1(\_142_[4] ),
    .S(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__clkbuf_1 _12086_ (.A(_06069_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _12087_ (.A0(\_140_[5] ),
    .A1(\_142_[5] ),
    .S(_06068_),
    .X(_06070_));
 sky130_fd_sc_hd__clkbuf_1 _12088_ (.A(_06070_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _12089_ (.A0(\_140_[6] ),
    .A1(\_142_[6] ),
    .S(_06068_),
    .X(_06071_));
 sky130_fd_sc_hd__clkbuf_1 _12090_ (.A(_06071_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _12091_ (.A0(\_140_[7] ),
    .A1(\_142_[7] ),
    .S(_06068_),
    .X(_06072_));
 sky130_fd_sc_hd__clkbuf_1 _12092_ (.A(_06072_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _12093_ (.A0(\_140_[8] ),
    .A1(\_142_[8] ),
    .S(_06068_),
    .X(_06073_));
 sky130_fd_sc_hd__clkbuf_1 _12094_ (.A(_06073_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _12095_ (.A0(\_140_[9] ),
    .A1(\_142_[9] ),
    .S(_06068_),
    .X(_06074_));
 sky130_fd_sc_hd__clkbuf_1 _12096_ (.A(_06074_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _12097_ (.A0(\_140_[10] ),
    .A1(\_142_[10] ),
    .S(_06068_),
    .X(_06075_));
 sky130_fd_sc_hd__clkbuf_1 _12098_ (.A(_06075_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _12099_ (.A0(\_140_[11] ),
    .A1(\_142_[11] ),
    .S(_06068_),
    .X(_06076_));
 sky130_fd_sc_hd__clkbuf_1 _12100_ (.A(_06076_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _12101_ (.A0(\_140_[12] ),
    .A1(\_142_[12] ),
    .S(_06068_),
    .X(_06077_));
 sky130_fd_sc_hd__clkbuf_1 _12102_ (.A(_06077_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _12103_ (.A0(\_140_[13] ),
    .A1(\_142_[13] ),
    .S(_06068_),
    .X(_06078_));
 sky130_fd_sc_hd__clkbuf_1 _12104_ (.A(_06078_),
    .X(_00832_));
 sky130_fd_sc_hd__clkbuf_4 _12105_ (.A(_06004_),
    .X(_06079_));
 sky130_fd_sc_hd__mux2_1 _12106_ (.A0(\_140_[14] ),
    .A1(\_142_[14] ),
    .S(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__clkbuf_1 _12107_ (.A(_06080_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _12108_ (.A0(\_140_[15] ),
    .A1(\_142_[15] ),
    .S(_06079_),
    .X(_06081_));
 sky130_fd_sc_hd__clkbuf_1 _12109_ (.A(_06081_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _12110_ (.A0(\_140_[16] ),
    .A1(\_142_[16] ),
    .S(_06079_),
    .X(_06082_));
 sky130_fd_sc_hd__clkbuf_1 _12111_ (.A(_06082_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _12112_ (.A0(\_140_[17] ),
    .A1(\_142_[17] ),
    .S(_06079_),
    .X(_06083_));
 sky130_fd_sc_hd__clkbuf_1 _12113_ (.A(_06083_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _12114_ (.A0(\_140_[18] ),
    .A1(\_142_[18] ),
    .S(_06079_),
    .X(_06084_));
 sky130_fd_sc_hd__clkbuf_1 _12115_ (.A(_06084_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _12116_ (.A0(\_140_[19] ),
    .A1(\_142_[19] ),
    .S(_06079_),
    .X(_06085_));
 sky130_fd_sc_hd__clkbuf_1 _12117_ (.A(_06085_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _12118_ (.A0(\_140_[20] ),
    .A1(\_142_[20] ),
    .S(_06079_),
    .X(_06086_));
 sky130_fd_sc_hd__clkbuf_1 _12119_ (.A(_06086_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _12120_ (.A0(\_140_[21] ),
    .A1(\_142_[21] ),
    .S(_06079_),
    .X(_06087_));
 sky130_fd_sc_hd__clkbuf_1 _12121_ (.A(_06087_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _12122_ (.A0(\_140_[22] ),
    .A1(\_142_[22] ),
    .S(_06079_),
    .X(_06088_));
 sky130_fd_sc_hd__clkbuf_1 _12123_ (.A(_06088_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _12124_ (.A0(\_140_[23] ),
    .A1(\_142_[23] ),
    .S(_06079_),
    .X(_06089_));
 sky130_fd_sc_hd__clkbuf_1 _12125_ (.A(_06089_),
    .X(_00842_));
 sky130_fd_sc_hd__buf_4 _12126_ (.A(_06004_),
    .X(_06090_));
 sky130_fd_sc_hd__mux2_1 _12127_ (.A0(\_140_[24] ),
    .A1(\_142_[24] ),
    .S(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__clkbuf_1 _12128_ (.A(_06091_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _12129_ (.A0(\_140_[25] ),
    .A1(\_142_[25] ),
    .S(_06090_),
    .X(_06092_));
 sky130_fd_sc_hd__clkbuf_1 _12130_ (.A(_06092_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _12131_ (.A0(\_140_[26] ),
    .A1(\_142_[26] ),
    .S(_06090_),
    .X(_06093_));
 sky130_fd_sc_hd__clkbuf_1 _12132_ (.A(_06093_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _12133_ (.A0(\_140_[27] ),
    .A1(\_142_[27] ),
    .S(_06090_),
    .X(_06094_));
 sky130_fd_sc_hd__clkbuf_1 _12134_ (.A(_06094_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _12135_ (.A0(\_140_[28] ),
    .A1(\_142_[28] ),
    .S(_06090_),
    .X(_06095_));
 sky130_fd_sc_hd__clkbuf_1 _12136_ (.A(_06095_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _12137_ (.A0(\_140_[29] ),
    .A1(\_142_[29] ),
    .S(_06090_),
    .X(_06096_));
 sky130_fd_sc_hd__clkbuf_1 _12138_ (.A(_06096_),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _12139_ (.A0(\_140_[30] ),
    .A1(\_142_[30] ),
    .S(_06090_),
    .X(_06097_));
 sky130_fd_sc_hd__clkbuf_1 _12140_ (.A(_06097_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _12141_ (.A0(\_140_[31] ),
    .A1(\_142_[31] ),
    .S(_06090_),
    .X(_06098_));
 sky130_fd_sc_hd__clkbuf_1 _12142_ (.A(_06098_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _12143_ (.A0(\_140_[0] ),
    .A1(\_138_[0] ),
    .S(_01394_),
    .X(_06099_));
 sky130_fd_sc_hd__clkbuf_1 _12144_ (.A(_06099_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _12145_ (.A0(\_140_[1] ),
    .A1(\_138_[1] ),
    .S(_01394_),
    .X(_06100_));
 sky130_fd_sc_hd__clkbuf_1 _12146_ (.A(_06100_),
    .X(_00852_));
 sky130_fd_sc_hd__clkbuf_4 _12147_ (.A(_01393_),
    .X(_06101_));
 sky130_fd_sc_hd__mux2_1 _12148_ (.A0(\_140_[2] ),
    .A1(\_138_[2] ),
    .S(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__clkbuf_1 _12149_ (.A(_06102_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _12150_ (.A0(\_140_[3] ),
    .A1(\_138_[3] ),
    .S(_06101_),
    .X(_06103_));
 sky130_fd_sc_hd__clkbuf_1 _12151_ (.A(_06103_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _12152_ (.A0(\_140_[4] ),
    .A1(\_138_[4] ),
    .S(_06101_),
    .X(_06104_));
 sky130_fd_sc_hd__clkbuf_1 _12153_ (.A(_06104_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _12154_ (.A0(\_140_[5] ),
    .A1(\_138_[5] ),
    .S(_06101_),
    .X(_06105_));
 sky130_fd_sc_hd__clkbuf_1 _12155_ (.A(_06105_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _12156_ (.A0(\_140_[6] ),
    .A1(\_138_[6] ),
    .S(_06101_),
    .X(_06106_));
 sky130_fd_sc_hd__clkbuf_1 _12157_ (.A(_06106_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _12158_ (.A0(\_140_[7] ),
    .A1(\_138_[7] ),
    .S(_06101_),
    .X(_06107_));
 sky130_fd_sc_hd__clkbuf_1 _12159_ (.A(_06107_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _12160_ (.A0(\_140_[8] ),
    .A1(\_138_[8] ),
    .S(_06101_),
    .X(_06108_));
 sky130_fd_sc_hd__clkbuf_1 _12161_ (.A(_06108_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _12162_ (.A0(\_140_[9] ),
    .A1(\_138_[9] ),
    .S(_06101_),
    .X(_06109_));
 sky130_fd_sc_hd__clkbuf_1 _12163_ (.A(_06109_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _12164_ (.A0(\_140_[10] ),
    .A1(\_138_[10] ),
    .S(_06101_),
    .X(_06110_));
 sky130_fd_sc_hd__clkbuf_1 _12165_ (.A(_06110_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _12166_ (.A0(\_140_[11] ),
    .A1(\_138_[11] ),
    .S(_06101_),
    .X(_06111_));
 sky130_fd_sc_hd__clkbuf_1 _12167_ (.A(_06111_),
    .X(_00862_));
 sky130_fd_sc_hd__clkbuf_4 _12168_ (.A(_01393_),
    .X(_06112_));
 sky130_fd_sc_hd__mux2_1 _12169_ (.A0(\_140_[12] ),
    .A1(\_138_[12] ),
    .S(_06112_),
    .X(_06113_));
 sky130_fd_sc_hd__clkbuf_1 _12170_ (.A(_06113_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _12171_ (.A0(\_140_[13] ),
    .A1(\_138_[13] ),
    .S(_06112_),
    .X(_06114_));
 sky130_fd_sc_hd__clkbuf_1 _12172_ (.A(_06114_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(\_140_[14] ),
    .A1(\_138_[14] ),
    .S(_06112_),
    .X(_06115_));
 sky130_fd_sc_hd__clkbuf_1 _12174_ (.A(_06115_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(\_140_[15] ),
    .A1(\_138_[15] ),
    .S(_06112_),
    .X(_06116_));
 sky130_fd_sc_hd__clkbuf_1 _12176_ (.A(_06116_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _12177_ (.A0(\_140_[16] ),
    .A1(\_138_[16] ),
    .S(_06112_),
    .X(_06117_));
 sky130_fd_sc_hd__clkbuf_1 _12178_ (.A(_06117_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _12179_ (.A0(\_140_[17] ),
    .A1(\_138_[17] ),
    .S(_06112_),
    .X(_06118_));
 sky130_fd_sc_hd__clkbuf_1 _12180_ (.A(_06118_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _12181_ (.A0(\_140_[18] ),
    .A1(\_138_[18] ),
    .S(_06112_),
    .X(_06119_));
 sky130_fd_sc_hd__clkbuf_1 _12182_ (.A(_06119_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _12183_ (.A0(\_140_[19] ),
    .A1(\_138_[19] ),
    .S(_06112_),
    .X(_06120_));
 sky130_fd_sc_hd__clkbuf_1 _12184_ (.A(_06120_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _12185_ (.A0(\_140_[20] ),
    .A1(\_138_[20] ),
    .S(_06112_),
    .X(_06121_));
 sky130_fd_sc_hd__clkbuf_1 _12186_ (.A(_06121_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _12187_ (.A0(\_140_[21] ),
    .A1(\_138_[21] ),
    .S(_06112_),
    .X(_06122_));
 sky130_fd_sc_hd__clkbuf_1 _12188_ (.A(_06122_),
    .X(_00872_));
 sky130_fd_sc_hd__clkbuf_4 _12189_ (.A(_01393_),
    .X(_06123_));
 sky130_fd_sc_hd__mux2_1 _12190_ (.A0(\_140_[22] ),
    .A1(\_138_[22] ),
    .S(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__clkbuf_1 _12191_ (.A(_06124_),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _12192_ (.A0(\_140_[23] ),
    .A1(\_138_[23] ),
    .S(_06123_),
    .X(_06125_));
 sky130_fd_sc_hd__clkbuf_1 _12193_ (.A(_06125_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _12194_ (.A0(\_140_[24] ),
    .A1(\_138_[24] ),
    .S(_06123_),
    .X(_06126_));
 sky130_fd_sc_hd__clkbuf_1 _12195_ (.A(_06126_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _12196_ (.A0(\_140_[25] ),
    .A1(\_138_[25] ),
    .S(_06123_),
    .X(_06127_));
 sky130_fd_sc_hd__clkbuf_1 _12197_ (.A(_06127_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _12198_ (.A0(\_140_[26] ),
    .A1(\_138_[26] ),
    .S(_06123_),
    .X(_06128_));
 sky130_fd_sc_hd__clkbuf_1 _12199_ (.A(_06128_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _12200_ (.A0(\_140_[27] ),
    .A1(\_138_[27] ),
    .S(_06123_),
    .X(_06129_));
 sky130_fd_sc_hd__clkbuf_1 _12201_ (.A(_06129_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _12202_ (.A0(\_140_[28] ),
    .A1(\_138_[28] ),
    .S(_06123_),
    .X(_06130_));
 sky130_fd_sc_hd__clkbuf_1 _12203_ (.A(_06130_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _12204_ (.A0(\_140_[29] ),
    .A1(\_138_[29] ),
    .S(_06123_),
    .X(_06131_));
 sky130_fd_sc_hd__clkbuf_1 _12205_ (.A(_06131_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _12206_ (.A0(\_140_[30] ),
    .A1(\_138_[30] ),
    .S(_06123_),
    .X(_06132_));
 sky130_fd_sc_hd__clkbuf_1 _12207_ (.A(_06132_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _12208_ (.A0(\_140_[31] ),
    .A1(\_138_[31] ),
    .S(_06123_),
    .X(_06133_));
 sky130_fd_sc_hd__clkbuf_1 _12209_ (.A(_06133_),
    .X(_00882_));
 sky130_fd_sc_hd__clkbuf_4 _12210_ (.A(_01393_),
    .X(_06134_));
 sky130_fd_sc_hd__mux2_1 _12211_ (.A0(\_138_[0] ),
    .A1(\_136_[0] ),
    .S(_06134_),
    .X(_06135_));
 sky130_fd_sc_hd__clkbuf_1 _12212_ (.A(_06135_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _12213_ (.A0(\_138_[1] ),
    .A1(\_136_[1] ),
    .S(_06134_),
    .X(_06136_));
 sky130_fd_sc_hd__clkbuf_1 _12214_ (.A(_06136_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _12215_ (.A0(\_138_[2] ),
    .A1(\_136_[2] ),
    .S(_06134_),
    .X(_06137_));
 sky130_fd_sc_hd__clkbuf_1 _12216_ (.A(_06137_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _12217_ (.A0(\_138_[3] ),
    .A1(\_136_[3] ),
    .S(_06134_),
    .X(_06138_));
 sky130_fd_sc_hd__clkbuf_1 _12218_ (.A(_06138_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _12219_ (.A0(\_138_[4] ),
    .A1(\_136_[4] ),
    .S(_06134_),
    .X(_06139_));
 sky130_fd_sc_hd__clkbuf_1 _12220_ (.A(_06139_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _12221_ (.A0(\_138_[5] ),
    .A1(\_136_[5] ),
    .S(_06134_),
    .X(_06140_));
 sky130_fd_sc_hd__clkbuf_1 _12222_ (.A(_06140_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _12223_ (.A0(\_138_[6] ),
    .A1(\_136_[6] ),
    .S(_06134_),
    .X(_06141_));
 sky130_fd_sc_hd__clkbuf_1 _12224_ (.A(_06141_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _12225_ (.A0(\_138_[7] ),
    .A1(\_136_[7] ),
    .S(_06134_),
    .X(_06142_));
 sky130_fd_sc_hd__clkbuf_1 _12226_ (.A(_06142_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _12227_ (.A0(\_138_[8] ),
    .A1(\_136_[8] ),
    .S(_06134_),
    .X(_06143_));
 sky130_fd_sc_hd__clkbuf_1 _12228_ (.A(_06143_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _12229_ (.A0(\_138_[9] ),
    .A1(\_136_[9] ),
    .S(_06134_),
    .X(_06144_));
 sky130_fd_sc_hd__clkbuf_1 _12230_ (.A(_06144_),
    .X(_00892_));
 sky130_fd_sc_hd__clkbuf_4 _12231_ (.A(_01393_),
    .X(_06145_));
 sky130_fd_sc_hd__mux2_1 _12232_ (.A0(\_138_[10] ),
    .A1(\_136_[10] ),
    .S(_06145_),
    .X(_06146_));
 sky130_fd_sc_hd__clkbuf_1 _12233_ (.A(_06146_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _12234_ (.A0(\_138_[11] ),
    .A1(\_136_[11] ),
    .S(_06145_),
    .X(_06147_));
 sky130_fd_sc_hd__clkbuf_1 _12235_ (.A(_06147_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _12236_ (.A0(\_138_[12] ),
    .A1(\_136_[12] ),
    .S(_06145_),
    .X(_06148_));
 sky130_fd_sc_hd__clkbuf_1 _12237_ (.A(_06148_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _12238_ (.A0(\_138_[13] ),
    .A1(\_136_[13] ),
    .S(_06145_),
    .X(_06149_));
 sky130_fd_sc_hd__clkbuf_1 _12239_ (.A(_06149_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(\_138_[14] ),
    .A1(\_136_[14] ),
    .S(_06145_),
    .X(_06150_));
 sky130_fd_sc_hd__clkbuf_1 _12241_ (.A(_06150_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _12242_ (.A0(\_138_[15] ),
    .A1(\_136_[15] ),
    .S(_06145_),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_1 _12243_ (.A(_06151_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _12244_ (.A0(\_138_[16] ),
    .A1(\_136_[16] ),
    .S(_06145_),
    .X(_06152_));
 sky130_fd_sc_hd__clkbuf_1 _12245_ (.A(_06152_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _12246_ (.A0(\_138_[17] ),
    .A1(\_136_[17] ),
    .S(_06145_),
    .X(_06153_));
 sky130_fd_sc_hd__clkbuf_1 _12247_ (.A(_06153_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _12248_ (.A0(\_138_[18] ),
    .A1(\_136_[18] ),
    .S(_06145_),
    .X(_06154_));
 sky130_fd_sc_hd__clkbuf_1 _12249_ (.A(_06154_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _12250_ (.A0(\_138_[19] ),
    .A1(\_136_[19] ),
    .S(_06145_),
    .X(_06155_));
 sky130_fd_sc_hd__clkbuf_1 _12251_ (.A(_06155_),
    .X(_00902_));
 sky130_fd_sc_hd__clkbuf_4 _12252_ (.A(_01393_),
    .X(_06156_));
 sky130_fd_sc_hd__mux2_1 _12253_ (.A0(\_138_[20] ),
    .A1(\_136_[20] ),
    .S(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__clkbuf_1 _12254_ (.A(_06157_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _12255_ (.A0(\_138_[21] ),
    .A1(\_136_[21] ),
    .S(_06156_),
    .X(_06158_));
 sky130_fd_sc_hd__clkbuf_1 _12256_ (.A(_06158_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _12257_ (.A0(\_138_[22] ),
    .A1(\_136_[22] ),
    .S(_06156_),
    .X(_06159_));
 sky130_fd_sc_hd__clkbuf_1 _12258_ (.A(_06159_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _12259_ (.A0(\_138_[23] ),
    .A1(\_136_[23] ),
    .S(_06156_),
    .X(_06160_));
 sky130_fd_sc_hd__clkbuf_1 _12260_ (.A(_06160_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _12261_ (.A0(\_138_[24] ),
    .A1(\_136_[24] ),
    .S(_06156_),
    .X(_06161_));
 sky130_fd_sc_hd__clkbuf_1 _12262_ (.A(_06161_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _12263_ (.A0(\_138_[25] ),
    .A1(\_136_[25] ),
    .S(_06156_),
    .X(_06162_));
 sky130_fd_sc_hd__clkbuf_1 _12264_ (.A(_06162_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _12265_ (.A0(\_138_[26] ),
    .A1(\_136_[26] ),
    .S(_06156_),
    .X(_06163_));
 sky130_fd_sc_hd__clkbuf_1 _12266_ (.A(_06163_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _12267_ (.A0(\_138_[27] ),
    .A1(\_136_[27] ),
    .S(_06156_),
    .X(_06164_));
 sky130_fd_sc_hd__clkbuf_1 _12268_ (.A(_06164_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _12269_ (.A0(\_138_[28] ),
    .A1(\_136_[28] ),
    .S(_06156_),
    .X(_06165_));
 sky130_fd_sc_hd__clkbuf_1 _12270_ (.A(_06165_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _12271_ (.A0(\_138_[29] ),
    .A1(\_136_[29] ),
    .S(_06156_),
    .X(_06166_));
 sky130_fd_sc_hd__clkbuf_1 _12272_ (.A(_06166_),
    .X(_00912_));
 sky130_fd_sc_hd__clkbuf_4 _12273_ (.A(_01393_),
    .X(_06167_));
 sky130_fd_sc_hd__mux2_1 _12274_ (.A0(\_138_[30] ),
    .A1(\_136_[30] ),
    .S(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__clkbuf_1 _12275_ (.A(_06168_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _12276_ (.A0(\_138_[31] ),
    .A1(\_136_[31] ),
    .S(_06167_),
    .X(_06169_));
 sky130_fd_sc_hd__clkbuf_1 _12277_ (.A(_06169_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _12278_ (.A0(\_136_[0] ),
    .A1(\_134_[0] ),
    .S(_06167_),
    .X(_06170_));
 sky130_fd_sc_hd__clkbuf_1 _12279_ (.A(_06170_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _12280_ (.A0(\_136_[1] ),
    .A1(\_134_[1] ),
    .S(_06167_),
    .X(_06171_));
 sky130_fd_sc_hd__clkbuf_1 _12281_ (.A(_06171_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _12282_ (.A0(\_136_[2] ),
    .A1(\_134_[2] ),
    .S(_06167_),
    .X(_06172_));
 sky130_fd_sc_hd__clkbuf_1 _12283_ (.A(_06172_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _12284_ (.A0(\_136_[3] ),
    .A1(\_134_[3] ),
    .S(_06167_),
    .X(_06173_));
 sky130_fd_sc_hd__clkbuf_1 _12285_ (.A(_06173_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _12286_ (.A0(\_136_[4] ),
    .A1(\_134_[4] ),
    .S(_06167_),
    .X(_06174_));
 sky130_fd_sc_hd__clkbuf_1 _12287_ (.A(_06174_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _12288_ (.A0(\_136_[5] ),
    .A1(\_134_[5] ),
    .S(_06167_),
    .X(_06175_));
 sky130_fd_sc_hd__clkbuf_1 _12289_ (.A(_06175_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _12290_ (.A0(\_136_[6] ),
    .A1(\_134_[6] ),
    .S(_06167_),
    .X(_06176_));
 sky130_fd_sc_hd__clkbuf_1 _12291_ (.A(_06176_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _12292_ (.A0(\_136_[7] ),
    .A1(\_134_[7] ),
    .S(_06167_),
    .X(_06177_));
 sky130_fd_sc_hd__clkbuf_1 _12293_ (.A(_06177_),
    .X(_00922_));
 sky130_fd_sc_hd__buf_4 _12294_ (.A(_01393_),
    .X(_06178_));
 sky130_fd_sc_hd__mux2_1 _12295_ (.A0(\_136_[8] ),
    .A1(\_134_[8] ),
    .S(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__clkbuf_1 _12296_ (.A(_06179_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _12297_ (.A0(\_136_[9] ),
    .A1(\_134_[9] ),
    .S(_06178_),
    .X(_06180_));
 sky130_fd_sc_hd__clkbuf_1 _12298_ (.A(_06180_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _12299_ (.A0(\_136_[10] ),
    .A1(\_134_[10] ),
    .S(_06178_),
    .X(_06181_));
 sky130_fd_sc_hd__clkbuf_1 _12300_ (.A(_06181_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _12301_ (.A0(\_136_[11] ),
    .A1(\_134_[11] ),
    .S(_06178_),
    .X(_06182_));
 sky130_fd_sc_hd__clkbuf_1 _12302_ (.A(_06182_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _12303_ (.A0(\_136_[12] ),
    .A1(\_134_[12] ),
    .S(_06178_),
    .X(_06183_));
 sky130_fd_sc_hd__clkbuf_1 _12304_ (.A(_06183_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _12305_ (.A0(\_136_[13] ),
    .A1(\_134_[13] ),
    .S(_06178_),
    .X(_06184_));
 sky130_fd_sc_hd__clkbuf_1 _12306_ (.A(_06184_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _12307_ (.A0(\_136_[14] ),
    .A1(\_134_[14] ),
    .S(_06178_),
    .X(_06185_));
 sky130_fd_sc_hd__clkbuf_1 _12308_ (.A(_06185_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _12309_ (.A0(\_136_[15] ),
    .A1(\_134_[15] ),
    .S(_06178_),
    .X(_06186_));
 sky130_fd_sc_hd__clkbuf_1 _12310_ (.A(_06186_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _12311_ (.A0(\_136_[16] ),
    .A1(\_134_[16] ),
    .S(_06178_),
    .X(_06187_));
 sky130_fd_sc_hd__clkbuf_1 _12312_ (.A(_06187_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _12313_ (.A0(\_136_[17] ),
    .A1(\_134_[17] ),
    .S(_06178_),
    .X(_06188_));
 sky130_fd_sc_hd__clkbuf_1 _12314_ (.A(_06188_),
    .X(_00932_));
 sky130_fd_sc_hd__clkbuf_4 _12315_ (.A(_01393_),
    .X(_06189_));
 sky130_fd_sc_hd__mux2_1 _12316_ (.A0(\_136_[18] ),
    .A1(\_134_[18] ),
    .S(_06189_),
    .X(_06190_));
 sky130_fd_sc_hd__clkbuf_1 _12317_ (.A(_06190_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _12318_ (.A0(\_136_[19] ),
    .A1(\_134_[19] ),
    .S(_06189_),
    .X(_06191_));
 sky130_fd_sc_hd__clkbuf_1 _12319_ (.A(_06191_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _12320_ (.A0(\_136_[20] ),
    .A1(\_134_[20] ),
    .S(_06189_),
    .X(_06192_));
 sky130_fd_sc_hd__clkbuf_1 _12321_ (.A(_06192_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _12322_ (.A0(\_136_[21] ),
    .A1(\_134_[21] ),
    .S(_06189_),
    .X(_06193_));
 sky130_fd_sc_hd__clkbuf_1 _12323_ (.A(_06193_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _12324_ (.A0(\_136_[22] ),
    .A1(\_134_[22] ),
    .S(_06189_),
    .X(_06194_));
 sky130_fd_sc_hd__clkbuf_1 _12325_ (.A(_06194_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _12326_ (.A0(\_136_[23] ),
    .A1(\_134_[23] ),
    .S(_06189_),
    .X(_06195_));
 sky130_fd_sc_hd__clkbuf_1 _12327_ (.A(_06195_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _12328_ (.A0(\_136_[24] ),
    .A1(\_134_[24] ),
    .S(_06189_),
    .X(_06196_));
 sky130_fd_sc_hd__clkbuf_1 _12329_ (.A(_06196_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _12330_ (.A0(\_136_[25] ),
    .A1(\_134_[25] ),
    .S(_06189_),
    .X(_06197_));
 sky130_fd_sc_hd__clkbuf_1 _12331_ (.A(_06197_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _12332_ (.A0(\_136_[26] ),
    .A1(\_134_[26] ),
    .S(_06189_),
    .X(_06198_));
 sky130_fd_sc_hd__clkbuf_1 _12333_ (.A(_06198_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _12334_ (.A0(\_136_[27] ),
    .A1(\_134_[27] ),
    .S(_06189_),
    .X(_06199_));
 sky130_fd_sc_hd__clkbuf_1 _12335_ (.A(_06199_),
    .X(_00942_));
 sky130_fd_sc_hd__buf_4 _12336_ (.A(_01366_),
    .X(_06200_));
 sky130_fd_sc_hd__clkbuf_4 _12337_ (.A(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__mux2_1 _12338_ (.A0(\_136_[28] ),
    .A1(\_134_[28] ),
    .S(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__clkbuf_1 _12339_ (.A(_06202_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _12340_ (.A0(\_136_[29] ),
    .A1(\_134_[29] ),
    .S(_06201_),
    .X(_06203_));
 sky130_fd_sc_hd__clkbuf_1 _12341_ (.A(_06203_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _12342_ (.A0(\_136_[30] ),
    .A1(\_134_[30] ),
    .S(_06201_),
    .X(_06204_));
 sky130_fd_sc_hd__clkbuf_1 _12343_ (.A(_06204_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _12344_ (.A0(\_136_[31] ),
    .A1(\_134_[31] ),
    .S(_06201_),
    .X(_06205_));
 sky130_fd_sc_hd__clkbuf_1 _12345_ (.A(_06205_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _12346_ (.A0(\_132_[0] ),
    .A1(\_134_[0] ),
    .S(_06090_),
    .X(_06206_));
 sky130_fd_sc_hd__clkbuf_1 _12347_ (.A(_06206_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _12348_ (.A0(\_132_[1] ),
    .A1(\_134_[1] ),
    .S(_06090_),
    .X(_06207_));
 sky130_fd_sc_hd__clkbuf_1 _12349_ (.A(_06207_),
    .X(_00948_));
 sky130_fd_sc_hd__buf_4 _12350_ (.A(_06004_),
    .X(_06208_));
 sky130_fd_sc_hd__mux2_1 _12351_ (.A0(\_132_[2] ),
    .A1(\_134_[2] ),
    .S(_06208_),
    .X(_06209_));
 sky130_fd_sc_hd__clkbuf_1 _12352_ (.A(_06209_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _12353_ (.A0(\_132_[3] ),
    .A1(\_134_[3] ),
    .S(_06208_),
    .X(_06210_));
 sky130_fd_sc_hd__clkbuf_1 _12354_ (.A(_06210_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _12355_ (.A0(\_132_[4] ),
    .A1(\_134_[4] ),
    .S(_06208_),
    .X(_06211_));
 sky130_fd_sc_hd__clkbuf_1 _12356_ (.A(_06211_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _12357_ (.A0(\_132_[5] ),
    .A1(\_134_[5] ),
    .S(_06208_),
    .X(_06212_));
 sky130_fd_sc_hd__clkbuf_1 _12358_ (.A(_06212_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _12359_ (.A0(\_132_[6] ),
    .A1(\_134_[6] ),
    .S(_06208_),
    .X(_06213_));
 sky130_fd_sc_hd__clkbuf_1 _12360_ (.A(_06213_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _12361_ (.A0(\_132_[7] ),
    .A1(\_134_[7] ),
    .S(_06208_),
    .X(_06214_));
 sky130_fd_sc_hd__clkbuf_1 _12362_ (.A(_06214_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _12363_ (.A0(\_132_[8] ),
    .A1(\_134_[8] ),
    .S(_06208_),
    .X(_06215_));
 sky130_fd_sc_hd__clkbuf_1 _12364_ (.A(_06215_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _12365_ (.A0(\_132_[9] ),
    .A1(\_134_[9] ),
    .S(_06208_),
    .X(_06216_));
 sky130_fd_sc_hd__clkbuf_1 _12366_ (.A(_06216_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _12367_ (.A0(\_132_[10] ),
    .A1(\_134_[10] ),
    .S(_06208_),
    .X(_06217_));
 sky130_fd_sc_hd__clkbuf_1 _12368_ (.A(_06217_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _12369_ (.A0(\_132_[11] ),
    .A1(\_134_[11] ),
    .S(_06208_),
    .X(_06218_));
 sky130_fd_sc_hd__clkbuf_1 _12370_ (.A(_06218_),
    .X(_00958_));
 sky130_fd_sc_hd__clkbuf_4 _12371_ (.A(_06004_),
    .X(_06219_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(\_132_[12] ),
    .A1(\_134_[12] ),
    .S(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__clkbuf_1 _12373_ (.A(_06220_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _12374_ (.A0(\_132_[13] ),
    .A1(\_134_[13] ),
    .S(_06219_),
    .X(_06221_));
 sky130_fd_sc_hd__clkbuf_1 _12375_ (.A(_06221_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _12376_ (.A0(\_132_[14] ),
    .A1(\_134_[14] ),
    .S(_06219_),
    .X(_06222_));
 sky130_fd_sc_hd__clkbuf_1 _12377_ (.A(_06222_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(\_132_[15] ),
    .A1(\_134_[15] ),
    .S(_06219_),
    .X(_06223_));
 sky130_fd_sc_hd__clkbuf_1 _12379_ (.A(_06223_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(\_132_[16] ),
    .A1(\_134_[16] ),
    .S(_06219_),
    .X(_06224_));
 sky130_fd_sc_hd__clkbuf_1 _12381_ (.A(_06224_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(\_132_[17] ),
    .A1(\_134_[17] ),
    .S(_06219_),
    .X(_06225_));
 sky130_fd_sc_hd__clkbuf_1 _12383_ (.A(_06225_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(\_132_[18] ),
    .A1(\_134_[18] ),
    .S(_06219_),
    .X(_06226_));
 sky130_fd_sc_hd__clkbuf_1 _12385_ (.A(_06226_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _12386_ (.A0(\_132_[19] ),
    .A1(\_134_[19] ),
    .S(_06219_),
    .X(_06227_));
 sky130_fd_sc_hd__clkbuf_1 _12387_ (.A(_06227_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(\_132_[20] ),
    .A1(\_134_[20] ),
    .S(_06219_),
    .X(_06228_));
 sky130_fd_sc_hd__clkbuf_1 _12389_ (.A(_06228_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(\_132_[21] ),
    .A1(\_134_[21] ),
    .S(_06219_),
    .X(_06229_));
 sky130_fd_sc_hd__clkbuf_1 _12391_ (.A(_06229_),
    .X(_00968_));
 sky130_fd_sc_hd__clkbuf_4 _12392_ (.A(_06004_),
    .X(_06230_));
 sky130_fd_sc_hd__mux2_1 _12393_ (.A0(\_132_[22] ),
    .A1(\_134_[22] ),
    .S(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__clkbuf_1 _12394_ (.A(_06231_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _12395_ (.A0(\_132_[23] ),
    .A1(\_134_[23] ),
    .S(_06230_),
    .X(_06232_));
 sky130_fd_sc_hd__clkbuf_1 _12396_ (.A(_06232_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _12397_ (.A0(\_132_[24] ),
    .A1(\_134_[24] ),
    .S(_06230_),
    .X(_06233_));
 sky130_fd_sc_hd__clkbuf_1 _12398_ (.A(_06233_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _12399_ (.A0(\_132_[25] ),
    .A1(\_134_[25] ),
    .S(_06230_),
    .X(_06234_));
 sky130_fd_sc_hd__clkbuf_1 _12400_ (.A(_06234_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _12401_ (.A0(\_132_[26] ),
    .A1(\_134_[26] ),
    .S(_06230_),
    .X(_06235_));
 sky130_fd_sc_hd__clkbuf_1 _12402_ (.A(_06235_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _12403_ (.A0(\_132_[27] ),
    .A1(\_134_[27] ),
    .S(_06230_),
    .X(_06236_));
 sky130_fd_sc_hd__clkbuf_1 _12404_ (.A(_06236_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _12405_ (.A0(\_132_[28] ),
    .A1(\_134_[28] ),
    .S(_06230_),
    .X(_06237_));
 sky130_fd_sc_hd__clkbuf_1 _12406_ (.A(_06237_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _12407_ (.A0(\_132_[29] ),
    .A1(\_134_[29] ),
    .S(_06230_),
    .X(_06238_));
 sky130_fd_sc_hd__clkbuf_1 _12408_ (.A(_06238_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _12409_ (.A0(\_132_[30] ),
    .A1(\_134_[30] ),
    .S(_06230_),
    .X(_06239_));
 sky130_fd_sc_hd__clkbuf_1 _12410_ (.A(_06239_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _12411_ (.A0(\_132_[31] ),
    .A1(\_134_[31] ),
    .S(_06230_),
    .X(_06240_));
 sky130_fd_sc_hd__clkbuf_1 _12412_ (.A(_06240_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _12413_ (.A0(\_132_[0] ),
    .A1(\_130_[0] ),
    .S(_06201_),
    .X(_06241_));
 sky130_fd_sc_hd__clkbuf_1 _12414_ (.A(_06241_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _12415_ (.A0(\_132_[1] ),
    .A1(\_130_[1] ),
    .S(_06201_),
    .X(_06242_));
 sky130_fd_sc_hd__clkbuf_1 _12416_ (.A(_06242_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _12417_ (.A0(\_132_[2] ),
    .A1(\_130_[2] ),
    .S(_06201_),
    .X(_06243_));
 sky130_fd_sc_hd__clkbuf_1 _12418_ (.A(_06243_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _12419_ (.A0(\_132_[3] ),
    .A1(\_130_[3] ),
    .S(_06201_),
    .X(_06244_));
 sky130_fd_sc_hd__clkbuf_1 _12420_ (.A(_06244_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _12421_ (.A0(\_132_[4] ),
    .A1(\_130_[4] ),
    .S(_06201_),
    .X(_06245_));
 sky130_fd_sc_hd__clkbuf_1 _12422_ (.A(_06245_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _12423_ (.A0(\_132_[5] ),
    .A1(\_130_[5] ),
    .S(_06201_),
    .X(_06246_));
 sky130_fd_sc_hd__clkbuf_1 _12424_ (.A(_06246_),
    .X(_00984_));
 sky130_fd_sc_hd__clkbuf_8 _12425_ (.A(_06200_),
    .X(_06247_));
 sky130_fd_sc_hd__mux2_1 _12426_ (.A0(\_132_[6] ),
    .A1(\_130_[6] ),
    .S(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__clkbuf_1 _12427_ (.A(_06248_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _12428_ (.A0(\_132_[7] ),
    .A1(\_130_[7] ),
    .S(_06247_),
    .X(_06249_));
 sky130_fd_sc_hd__clkbuf_1 _12429_ (.A(_06249_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _12430_ (.A0(\_132_[8] ),
    .A1(\_130_[8] ),
    .S(_06247_),
    .X(_06250_));
 sky130_fd_sc_hd__clkbuf_1 _12431_ (.A(_06250_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _12432_ (.A0(\_132_[9] ),
    .A1(\_130_[9] ),
    .S(_06247_),
    .X(_06251_));
 sky130_fd_sc_hd__clkbuf_1 _12433_ (.A(_06251_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _12434_ (.A0(\_132_[10] ),
    .A1(\_130_[10] ),
    .S(_06247_),
    .X(_06252_));
 sky130_fd_sc_hd__clkbuf_1 _12435_ (.A(_06252_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _12436_ (.A0(\_132_[11] ),
    .A1(\_130_[11] ),
    .S(_06247_),
    .X(_06253_));
 sky130_fd_sc_hd__clkbuf_1 _12437_ (.A(_06253_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _12438_ (.A0(\_132_[12] ),
    .A1(\_130_[12] ),
    .S(_06247_),
    .X(_06254_));
 sky130_fd_sc_hd__clkbuf_1 _12439_ (.A(_06254_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _12440_ (.A0(\_132_[13] ),
    .A1(\_130_[13] ),
    .S(_06247_),
    .X(_06255_));
 sky130_fd_sc_hd__clkbuf_1 _12441_ (.A(_06255_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _12442_ (.A0(\_132_[14] ),
    .A1(\_130_[14] ),
    .S(_06247_),
    .X(_06256_));
 sky130_fd_sc_hd__clkbuf_1 _12443_ (.A(_06256_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _12444_ (.A0(\_132_[15] ),
    .A1(\_130_[15] ),
    .S(_06247_),
    .X(_06257_));
 sky130_fd_sc_hd__clkbuf_1 _12445_ (.A(_06257_),
    .X(_00994_));
 sky130_fd_sc_hd__buf_4 _12446_ (.A(_06200_),
    .X(_06258_));
 sky130_fd_sc_hd__mux2_1 _12447_ (.A0(\_132_[16] ),
    .A1(\_130_[16] ),
    .S(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__clkbuf_1 _12448_ (.A(_06259_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _12449_ (.A0(\_132_[17] ),
    .A1(\_130_[17] ),
    .S(_06258_),
    .X(_06260_));
 sky130_fd_sc_hd__clkbuf_1 _12450_ (.A(_06260_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(\_132_[18] ),
    .A1(\_130_[18] ),
    .S(_06258_),
    .X(_06261_));
 sky130_fd_sc_hd__clkbuf_1 _12452_ (.A(_06261_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _12453_ (.A0(\_132_[19] ),
    .A1(\_130_[19] ),
    .S(_06258_),
    .X(_06262_));
 sky130_fd_sc_hd__clkbuf_1 _12454_ (.A(_06262_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(\_132_[20] ),
    .A1(\_130_[20] ),
    .S(_06258_),
    .X(_06263_));
 sky130_fd_sc_hd__clkbuf_1 _12456_ (.A(_06263_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _12457_ (.A0(\_132_[21] ),
    .A1(\_130_[21] ),
    .S(_06258_),
    .X(_06264_));
 sky130_fd_sc_hd__clkbuf_1 _12458_ (.A(_06264_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _12459_ (.A0(\_132_[22] ),
    .A1(\_130_[22] ),
    .S(_06258_),
    .X(_06265_));
 sky130_fd_sc_hd__clkbuf_1 _12460_ (.A(_06265_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _12461_ (.A0(\_132_[23] ),
    .A1(\_130_[23] ),
    .S(_06258_),
    .X(_06266_));
 sky130_fd_sc_hd__clkbuf_1 _12462_ (.A(_06266_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _12463_ (.A0(\_132_[24] ),
    .A1(\_130_[24] ),
    .S(_06258_),
    .X(_06267_));
 sky130_fd_sc_hd__clkbuf_1 _12464_ (.A(_06267_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _12465_ (.A0(\_132_[25] ),
    .A1(\_130_[25] ),
    .S(_06258_),
    .X(_06268_));
 sky130_fd_sc_hd__clkbuf_1 _12466_ (.A(_06268_),
    .X(_01004_));
 sky130_fd_sc_hd__clkbuf_4 _12467_ (.A(_06200_),
    .X(_06269_));
 sky130_fd_sc_hd__mux2_1 _12468_ (.A0(\_132_[26] ),
    .A1(\_130_[26] ),
    .S(_06269_),
    .X(_06270_));
 sky130_fd_sc_hd__clkbuf_1 _12469_ (.A(_06270_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _12470_ (.A0(\_132_[27] ),
    .A1(\_130_[27] ),
    .S(_06269_),
    .X(_06271_));
 sky130_fd_sc_hd__clkbuf_1 _12471_ (.A(_06271_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(\_132_[28] ),
    .A1(\_130_[28] ),
    .S(_06269_),
    .X(_06272_));
 sky130_fd_sc_hd__clkbuf_1 _12473_ (.A(_06272_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _12474_ (.A0(\_132_[29] ),
    .A1(\_130_[29] ),
    .S(_06269_),
    .X(_06273_));
 sky130_fd_sc_hd__clkbuf_1 _12475_ (.A(_06273_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(\_132_[30] ),
    .A1(\_130_[30] ),
    .S(_06269_),
    .X(_06274_));
 sky130_fd_sc_hd__clkbuf_1 _12477_ (.A(_06274_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _12478_ (.A0(\_132_[31] ),
    .A1(\_130_[31] ),
    .S(_06269_),
    .X(_06275_));
 sky130_fd_sc_hd__clkbuf_1 _12479_ (.A(_06275_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _12480_ (.A0(\_130_[0] ),
    .A1(\_128_[0] ),
    .S(_06269_),
    .X(_06276_));
 sky130_fd_sc_hd__clkbuf_1 _12481_ (.A(_06276_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _12482_ (.A0(\_130_[1] ),
    .A1(\_128_[1] ),
    .S(_06269_),
    .X(_06277_));
 sky130_fd_sc_hd__clkbuf_1 _12483_ (.A(_06277_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _12484_ (.A0(\_130_[2] ),
    .A1(\_128_[2] ),
    .S(_06269_),
    .X(_06278_));
 sky130_fd_sc_hd__clkbuf_1 _12485_ (.A(_06278_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _12486_ (.A0(\_130_[3] ),
    .A1(\_128_[3] ),
    .S(_06269_),
    .X(_06279_));
 sky130_fd_sc_hd__clkbuf_1 _12487_ (.A(_06279_),
    .X(_01014_));
 sky130_fd_sc_hd__buf_6 _12488_ (.A(_06200_),
    .X(_06280_));
 sky130_fd_sc_hd__mux2_1 _12489_ (.A0(\_130_[4] ),
    .A1(\_128_[4] ),
    .S(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__clkbuf_1 _12490_ (.A(_06281_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _12491_ (.A0(\_130_[5] ),
    .A1(\_128_[5] ),
    .S(_06280_),
    .X(_06282_));
 sky130_fd_sc_hd__clkbuf_1 _12492_ (.A(_06282_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _12493_ (.A0(\_130_[6] ),
    .A1(\_128_[6] ),
    .S(_06280_),
    .X(_06283_));
 sky130_fd_sc_hd__clkbuf_1 _12494_ (.A(_06283_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _12495_ (.A0(\_130_[7] ),
    .A1(\_128_[7] ),
    .S(_06280_),
    .X(_06284_));
 sky130_fd_sc_hd__clkbuf_1 _12496_ (.A(_06284_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _12497_ (.A0(\_130_[8] ),
    .A1(\_128_[8] ),
    .S(_06280_),
    .X(_06285_));
 sky130_fd_sc_hd__clkbuf_1 _12498_ (.A(_06285_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(\_130_[9] ),
    .A1(\_128_[9] ),
    .S(_06280_),
    .X(_06286_));
 sky130_fd_sc_hd__clkbuf_1 _12500_ (.A(_06286_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _12501_ (.A0(\_130_[10] ),
    .A1(\_128_[10] ),
    .S(_06280_),
    .X(_06287_));
 sky130_fd_sc_hd__clkbuf_1 _12502_ (.A(_06287_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _12503_ (.A0(\_130_[11] ),
    .A1(\_128_[11] ),
    .S(_06280_),
    .X(_06288_));
 sky130_fd_sc_hd__clkbuf_1 _12504_ (.A(_06288_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _12505_ (.A0(\_130_[12] ),
    .A1(\_128_[12] ),
    .S(_06280_),
    .X(_06289_));
 sky130_fd_sc_hd__clkbuf_1 _12506_ (.A(_06289_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _12507_ (.A0(\_130_[13] ),
    .A1(\_128_[13] ),
    .S(_06280_),
    .X(_06290_));
 sky130_fd_sc_hd__clkbuf_1 _12508_ (.A(_06290_),
    .X(_01024_));
 sky130_fd_sc_hd__clkbuf_4 _12509_ (.A(_06200_),
    .X(_06291_));
 sky130_fd_sc_hd__mux2_1 _12510_ (.A0(\_130_[14] ),
    .A1(\_128_[14] ),
    .S(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__clkbuf_1 _12511_ (.A(_06292_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _12512_ (.A0(\_130_[15] ),
    .A1(\_128_[15] ),
    .S(_06291_),
    .X(_06293_));
 sky130_fd_sc_hd__clkbuf_1 _12513_ (.A(_06293_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _12514_ (.A0(\_130_[16] ),
    .A1(\_128_[16] ),
    .S(_06291_),
    .X(_06294_));
 sky130_fd_sc_hd__clkbuf_1 _12515_ (.A(_06294_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _12516_ (.A0(\_130_[17] ),
    .A1(\_128_[17] ),
    .S(_06291_),
    .X(_06295_));
 sky130_fd_sc_hd__clkbuf_1 _12517_ (.A(_06295_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _12518_ (.A0(\_130_[18] ),
    .A1(\_128_[18] ),
    .S(_06291_),
    .X(_06296_));
 sky130_fd_sc_hd__clkbuf_1 _12519_ (.A(_06296_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _12520_ (.A0(\_130_[19] ),
    .A1(\_128_[19] ),
    .S(_06291_),
    .X(_06297_));
 sky130_fd_sc_hd__clkbuf_1 _12521_ (.A(_06297_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _12522_ (.A0(\_130_[20] ),
    .A1(\_128_[20] ),
    .S(_06291_),
    .X(_06298_));
 sky130_fd_sc_hd__clkbuf_1 _12523_ (.A(_06298_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _12524_ (.A0(\_130_[21] ),
    .A1(\_128_[21] ),
    .S(_06291_),
    .X(_06299_));
 sky130_fd_sc_hd__clkbuf_1 _12525_ (.A(_06299_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _12526_ (.A0(\_130_[22] ),
    .A1(\_128_[22] ),
    .S(_06291_),
    .X(_06300_));
 sky130_fd_sc_hd__clkbuf_1 _12527_ (.A(_06300_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _12528_ (.A0(\_130_[23] ),
    .A1(\_128_[23] ),
    .S(_06291_),
    .X(_06301_));
 sky130_fd_sc_hd__clkbuf_1 _12529_ (.A(_06301_),
    .X(_01034_));
 sky130_fd_sc_hd__clkbuf_4 _12530_ (.A(_06200_),
    .X(_06302_));
 sky130_fd_sc_hd__mux2_1 _12531_ (.A0(\_130_[24] ),
    .A1(\_128_[24] ),
    .S(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__clkbuf_1 _12532_ (.A(_06303_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _12533_ (.A0(\_130_[25] ),
    .A1(\_128_[25] ),
    .S(_06302_),
    .X(_06304_));
 sky130_fd_sc_hd__clkbuf_1 _12534_ (.A(_06304_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _12535_ (.A0(\_130_[26] ),
    .A1(\_128_[26] ),
    .S(_06302_),
    .X(_06305_));
 sky130_fd_sc_hd__clkbuf_1 _12536_ (.A(_06305_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _12537_ (.A0(\_130_[27] ),
    .A1(\_128_[27] ),
    .S(_06302_),
    .X(_06306_));
 sky130_fd_sc_hd__clkbuf_1 _12538_ (.A(_06306_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(\_130_[28] ),
    .A1(\_128_[28] ),
    .S(_06302_),
    .X(_06307_));
 sky130_fd_sc_hd__clkbuf_1 _12540_ (.A(_06307_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(\_130_[29] ),
    .A1(\_128_[29] ),
    .S(_06302_),
    .X(_06308_));
 sky130_fd_sc_hd__clkbuf_1 _12542_ (.A(_06308_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _12543_ (.A0(\_130_[30] ),
    .A1(\_128_[30] ),
    .S(_06302_),
    .X(_06309_));
 sky130_fd_sc_hd__clkbuf_1 _12544_ (.A(_06309_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _12545_ (.A0(\_130_[31] ),
    .A1(\_128_[31] ),
    .S(_06302_),
    .X(_06310_));
 sky130_fd_sc_hd__clkbuf_1 _12546_ (.A(_06310_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _12547_ (.A0(\_128_[0] ),
    .A1(\_126_[0] ),
    .S(_06302_),
    .X(_06311_));
 sky130_fd_sc_hd__clkbuf_1 _12548_ (.A(_06311_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _12549_ (.A0(\_128_[1] ),
    .A1(\_126_[1] ),
    .S(_06302_),
    .X(_06312_));
 sky130_fd_sc_hd__clkbuf_1 _12550_ (.A(_06312_),
    .X(_01044_));
 sky130_fd_sc_hd__buf_4 _12551_ (.A(_06200_),
    .X(_06313_));
 sky130_fd_sc_hd__mux2_1 _12552_ (.A0(\_128_[2] ),
    .A1(\_126_[2] ),
    .S(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__clkbuf_1 _12553_ (.A(_06314_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _12554_ (.A0(\_128_[3] ),
    .A1(\_126_[3] ),
    .S(_06313_),
    .X(_06315_));
 sky130_fd_sc_hd__clkbuf_1 _12555_ (.A(_06315_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _12556_ (.A0(\_128_[4] ),
    .A1(\_126_[4] ),
    .S(_06313_),
    .X(_06316_));
 sky130_fd_sc_hd__clkbuf_1 _12557_ (.A(_06316_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _12558_ (.A0(\_128_[5] ),
    .A1(\_126_[5] ),
    .S(_06313_),
    .X(_06317_));
 sky130_fd_sc_hd__clkbuf_1 _12559_ (.A(_06317_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _12560_ (.A0(\_128_[6] ),
    .A1(\_126_[6] ),
    .S(_06313_),
    .X(_06318_));
 sky130_fd_sc_hd__clkbuf_1 _12561_ (.A(_06318_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _12562_ (.A0(\_128_[7] ),
    .A1(\_126_[7] ),
    .S(_06313_),
    .X(_06319_));
 sky130_fd_sc_hd__clkbuf_1 _12563_ (.A(_06319_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _12564_ (.A0(\_128_[8] ),
    .A1(\_126_[8] ),
    .S(_06313_),
    .X(_06320_));
 sky130_fd_sc_hd__clkbuf_1 _12565_ (.A(_06320_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _12566_ (.A0(\_128_[9] ),
    .A1(\_126_[9] ),
    .S(_06313_),
    .X(_06321_));
 sky130_fd_sc_hd__clkbuf_1 _12567_ (.A(_06321_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _12568_ (.A0(\_128_[10] ),
    .A1(\_126_[10] ),
    .S(_06313_),
    .X(_06322_));
 sky130_fd_sc_hd__clkbuf_1 _12569_ (.A(_06322_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _12570_ (.A0(\_128_[11] ),
    .A1(\_126_[11] ),
    .S(_06313_),
    .X(_06323_));
 sky130_fd_sc_hd__clkbuf_1 _12571_ (.A(_06323_),
    .X(_01054_));
 sky130_fd_sc_hd__clkbuf_4 _12572_ (.A(_06200_),
    .X(_06324_));
 sky130_fd_sc_hd__mux2_1 _12573_ (.A0(\_128_[12] ),
    .A1(\_126_[12] ),
    .S(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__clkbuf_1 _12574_ (.A(_06325_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _12575_ (.A0(\_128_[13] ),
    .A1(\_126_[13] ),
    .S(_06324_),
    .X(_06326_));
 sky130_fd_sc_hd__clkbuf_1 _12576_ (.A(_06326_),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _12577_ (.A0(\_128_[14] ),
    .A1(\_126_[14] ),
    .S(_06324_),
    .X(_06327_));
 sky130_fd_sc_hd__clkbuf_1 _12578_ (.A(_06327_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _12579_ (.A0(\_128_[15] ),
    .A1(\_126_[15] ),
    .S(_06324_),
    .X(_06328_));
 sky130_fd_sc_hd__clkbuf_1 _12580_ (.A(_06328_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _12581_ (.A0(\_128_[16] ),
    .A1(\_126_[16] ),
    .S(_06324_),
    .X(_06329_));
 sky130_fd_sc_hd__clkbuf_1 _12582_ (.A(_06329_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _12583_ (.A0(\_128_[17] ),
    .A1(\_126_[17] ),
    .S(_06324_),
    .X(_06330_));
 sky130_fd_sc_hd__clkbuf_1 _12584_ (.A(_06330_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _12585_ (.A0(\_128_[18] ),
    .A1(\_126_[18] ),
    .S(_06324_),
    .X(_06331_));
 sky130_fd_sc_hd__clkbuf_1 _12586_ (.A(_06331_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(\_128_[19] ),
    .A1(\_126_[19] ),
    .S(_06324_),
    .X(_06332_));
 sky130_fd_sc_hd__clkbuf_1 _12588_ (.A(_06332_),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _12589_ (.A0(\_128_[20] ),
    .A1(\_126_[20] ),
    .S(_06324_),
    .X(_06333_));
 sky130_fd_sc_hd__clkbuf_1 _12590_ (.A(_06333_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _12591_ (.A0(\_128_[21] ),
    .A1(\_126_[21] ),
    .S(_06324_),
    .X(_06334_));
 sky130_fd_sc_hd__clkbuf_1 _12592_ (.A(_06334_),
    .X(_01064_));
 sky130_fd_sc_hd__buf_4 _12593_ (.A(_06200_),
    .X(_06335_));
 sky130_fd_sc_hd__mux2_1 _12594_ (.A0(\_128_[22] ),
    .A1(\_126_[22] ),
    .S(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__clkbuf_1 _12595_ (.A(_06336_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(\_128_[23] ),
    .A1(\_126_[23] ),
    .S(_06335_),
    .X(_06337_));
 sky130_fd_sc_hd__clkbuf_1 _12597_ (.A(_06337_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _12598_ (.A0(\_128_[24] ),
    .A1(\_126_[24] ),
    .S(_06335_),
    .X(_06338_));
 sky130_fd_sc_hd__clkbuf_1 _12599_ (.A(_06338_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _12600_ (.A0(\_128_[25] ),
    .A1(\_126_[25] ),
    .S(_06335_),
    .X(_06339_));
 sky130_fd_sc_hd__clkbuf_1 _12601_ (.A(_06339_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _12602_ (.A0(\_128_[26] ),
    .A1(\_126_[26] ),
    .S(_06335_),
    .X(_06340_));
 sky130_fd_sc_hd__clkbuf_1 _12603_ (.A(_06340_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _12604_ (.A0(\_128_[27] ),
    .A1(\_126_[27] ),
    .S(_06335_),
    .X(_06341_));
 sky130_fd_sc_hd__clkbuf_1 _12605_ (.A(_06341_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _12606_ (.A0(\_128_[28] ),
    .A1(\_126_[28] ),
    .S(_06335_),
    .X(_06342_));
 sky130_fd_sc_hd__clkbuf_1 _12607_ (.A(_06342_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _12608_ (.A0(\_128_[29] ),
    .A1(\_126_[29] ),
    .S(_06335_),
    .X(_06343_));
 sky130_fd_sc_hd__clkbuf_1 _12609_ (.A(_06343_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _12610_ (.A0(\_128_[30] ),
    .A1(\_126_[30] ),
    .S(_06335_),
    .X(_06344_));
 sky130_fd_sc_hd__clkbuf_1 _12611_ (.A(_06344_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _12612_ (.A0(\_128_[31] ),
    .A1(\_126_[31] ),
    .S(_06335_),
    .X(_06345_));
 sky130_fd_sc_hd__clkbuf_1 _12613_ (.A(_06345_),
    .X(_01074_));
 sky130_fd_sc_hd__clkbuf_4 _12614_ (.A(_01392_),
    .X(_06346_));
 sky130_fd_sc_hd__mux2_1 _12615_ (.A0(\_126_[0] ),
    .A1(\_124_[0] ),
    .S(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__clkbuf_1 _12616_ (.A(_06347_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _12617_ (.A0(\_126_[1] ),
    .A1(\_124_[1] ),
    .S(_06346_),
    .X(_06348_));
 sky130_fd_sc_hd__clkbuf_1 _12618_ (.A(_06348_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _12619_ (.A0(\_126_[2] ),
    .A1(\_124_[2] ),
    .S(_06346_),
    .X(_06349_));
 sky130_fd_sc_hd__clkbuf_1 _12620_ (.A(_06349_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _12621_ (.A0(\_126_[3] ),
    .A1(\_124_[3] ),
    .S(_06346_),
    .X(_06350_));
 sky130_fd_sc_hd__clkbuf_1 _12622_ (.A(_06350_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _12623_ (.A0(\_126_[4] ),
    .A1(\_124_[4] ),
    .S(_06346_),
    .X(_06351_));
 sky130_fd_sc_hd__clkbuf_1 _12624_ (.A(_06351_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _12625_ (.A0(\_126_[5] ),
    .A1(\_124_[5] ),
    .S(_06346_),
    .X(_06352_));
 sky130_fd_sc_hd__clkbuf_1 _12626_ (.A(_06352_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _12627_ (.A0(\_126_[6] ),
    .A1(\_124_[6] ),
    .S(_06346_),
    .X(_06353_));
 sky130_fd_sc_hd__clkbuf_1 _12628_ (.A(_06353_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _12629_ (.A0(\_126_[7] ),
    .A1(\_124_[7] ),
    .S(_06346_),
    .X(_06354_));
 sky130_fd_sc_hd__clkbuf_1 _12630_ (.A(_06354_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _12631_ (.A0(\_126_[8] ),
    .A1(\_124_[8] ),
    .S(_06346_),
    .X(_06355_));
 sky130_fd_sc_hd__clkbuf_1 _12632_ (.A(_06355_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _12633_ (.A0(\_126_[9] ),
    .A1(\_124_[9] ),
    .S(_06346_),
    .X(_06356_));
 sky130_fd_sc_hd__clkbuf_1 _12634_ (.A(_06356_),
    .X(_01084_));
 sky130_fd_sc_hd__buf_4 _12635_ (.A(_01392_),
    .X(_06357_));
 sky130_fd_sc_hd__mux2_1 _12636_ (.A0(\_126_[10] ),
    .A1(\_124_[10] ),
    .S(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__clkbuf_1 _12637_ (.A(_06358_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _12638_ (.A0(\_126_[11] ),
    .A1(\_124_[11] ),
    .S(_06357_),
    .X(_06359_));
 sky130_fd_sc_hd__clkbuf_1 _12639_ (.A(_06359_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _12640_ (.A0(\_126_[12] ),
    .A1(\_124_[12] ),
    .S(_06357_),
    .X(_06360_));
 sky130_fd_sc_hd__clkbuf_1 _12641_ (.A(_06360_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _12642_ (.A0(\_126_[13] ),
    .A1(\_124_[13] ),
    .S(_06357_),
    .X(_06361_));
 sky130_fd_sc_hd__clkbuf_1 _12643_ (.A(_06361_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _12644_ (.A0(\_126_[14] ),
    .A1(\_124_[14] ),
    .S(_06357_),
    .X(_06362_));
 sky130_fd_sc_hd__clkbuf_1 _12645_ (.A(_06362_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _12646_ (.A0(\_126_[15] ),
    .A1(\_124_[15] ),
    .S(_06357_),
    .X(_06363_));
 sky130_fd_sc_hd__clkbuf_1 _12647_ (.A(_06363_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _12648_ (.A0(\_126_[16] ),
    .A1(\_124_[16] ),
    .S(_06357_),
    .X(_06364_));
 sky130_fd_sc_hd__clkbuf_1 _12649_ (.A(_06364_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _12650_ (.A0(\_126_[17] ),
    .A1(\_124_[17] ),
    .S(_06357_),
    .X(_06365_));
 sky130_fd_sc_hd__clkbuf_1 _12651_ (.A(_06365_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _12652_ (.A0(\_126_[18] ),
    .A1(\_124_[18] ),
    .S(_06357_),
    .X(_06366_));
 sky130_fd_sc_hd__clkbuf_1 _12653_ (.A(_06366_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _12654_ (.A0(\_126_[19] ),
    .A1(\_124_[19] ),
    .S(_06357_),
    .X(_06367_));
 sky130_fd_sc_hd__clkbuf_1 _12655_ (.A(_06367_),
    .X(_01094_));
 sky130_fd_sc_hd__buf_4 _12656_ (.A(_01392_),
    .X(_06368_));
 sky130_fd_sc_hd__mux2_1 _12657_ (.A0(\_126_[20] ),
    .A1(\_124_[20] ),
    .S(_06368_),
    .X(_06369_));
 sky130_fd_sc_hd__clkbuf_1 _12658_ (.A(_06369_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _12659_ (.A0(\_126_[21] ),
    .A1(\_124_[21] ),
    .S(_06368_),
    .X(_06370_));
 sky130_fd_sc_hd__clkbuf_1 _12660_ (.A(_06370_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _12661_ (.A0(\_126_[22] ),
    .A1(\_124_[22] ),
    .S(_06368_),
    .X(_06371_));
 sky130_fd_sc_hd__clkbuf_1 _12662_ (.A(_06371_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _12663_ (.A0(\_126_[23] ),
    .A1(\_124_[23] ),
    .S(_06368_),
    .X(_06372_));
 sky130_fd_sc_hd__clkbuf_1 _12664_ (.A(_06372_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _12665_ (.A0(\_126_[24] ),
    .A1(\_124_[24] ),
    .S(_06368_),
    .X(_06373_));
 sky130_fd_sc_hd__clkbuf_1 _12666_ (.A(_06373_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _12667_ (.A0(\_126_[25] ),
    .A1(\_124_[25] ),
    .S(_06368_),
    .X(_06374_));
 sky130_fd_sc_hd__clkbuf_1 _12668_ (.A(_06374_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _12669_ (.A0(\_126_[26] ),
    .A1(\_124_[26] ),
    .S(_06368_),
    .X(_06375_));
 sky130_fd_sc_hd__clkbuf_1 _12670_ (.A(_06375_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _12671_ (.A0(\_126_[27] ),
    .A1(\_124_[27] ),
    .S(_06368_),
    .X(_06376_));
 sky130_fd_sc_hd__clkbuf_1 _12672_ (.A(_06376_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _12673_ (.A0(\_126_[28] ),
    .A1(\_124_[28] ),
    .S(_06368_),
    .X(_06377_));
 sky130_fd_sc_hd__clkbuf_1 _12674_ (.A(_06377_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _12675_ (.A0(\_126_[29] ),
    .A1(\_124_[29] ),
    .S(_06368_),
    .X(_06378_));
 sky130_fd_sc_hd__clkbuf_1 _12676_ (.A(_06378_),
    .X(_01104_));
 sky130_fd_sc_hd__clkbuf_4 _12677_ (.A(_01392_),
    .X(_06379_));
 sky130_fd_sc_hd__mux2_1 _12678_ (.A0(\_126_[30] ),
    .A1(\_124_[30] ),
    .S(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__clkbuf_1 _12679_ (.A(_06380_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _12680_ (.A0(\_126_[31] ),
    .A1(\_124_[31] ),
    .S(_06379_),
    .X(_06381_));
 sky130_fd_sc_hd__clkbuf_1 _12681_ (.A(_06381_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _12682_ (.A0(\_124_[0] ),
    .A1(\_122_[0] ),
    .S(_06379_),
    .X(_06382_));
 sky130_fd_sc_hd__clkbuf_1 _12683_ (.A(_06382_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _12684_ (.A0(\_124_[1] ),
    .A1(\_122_[1] ),
    .S(_06379_),
    .X(_06383_));
 sky130_fd_sc_hd__clkbuf_1 _12685_ (.A(_06383_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _12686_ (.A0(\_124_[2] ),
    .A1(\_122_[2] ),
    .S(_06379_),
    .X(_06384_));
 sky130_fd_sc_hd__clkbuf_1 _12687_ (.A(_06384_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _12688_ (.A0(\_124_[3] ),
    .A1(\_122_[3] ),
    .S(_06379_),
    .X(_06385_));
 sky130_fd_sc_hd__clkbuf_1 _12689_ (.A(_06385_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _12690_ (.A0(\_124_[4] ),
    .A1(\_122_[4] ),
    .S(_06379_),
    .X(_06386_));
 sky130_fd_sc_hd__clkbuf_1 _12691_ (.A(_06386_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _12692_ (.A0(\_124_[5] ),
    .A1(\_122_[5] ),
    .S(_06379_),
    .X(_06387_));
 sky130_fd_sc_hd__clkbuf_1 _12693_ (.A(_06387_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _12694_ (.A0(\_124_[6] ),
    .A1(\_122_[6] ),
    .S(_06379_),
    .X(_06388_));
 sky130_fd_sc_hd__clkbuf_1 _12695_ (.A(_06388_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _12696_ (.A0(\_124_[7] ),
    .A1(\_122_[7] ),
    .S(_06379_),
    .X(_06389_));
 sky130_fd_sc_hd__clkbuf_1 _12697_ (.A(_06389_),
    .X(_01114_));
 sky130_fd_sc_hd__buf_6 _12698_ (.A(_01392_),
    .X(_06390_));
 sky130_fd_sc_hd__mux2_1 _12699_ (.A0(\_124_[8] ),
    .A1(\_122_[8] ),
    .S(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__clkbuf_1 _12700_ (.A(_06391_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _12701_ (.A0(\_124_[9] ),
    .A1(\_122_[9] ),
    .S(_06390_),
    .X(_06392_));
 sky130_fd_sc_hd__clkbuf_1 _12702_ (.A(_06392_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _12703_ (.A0(\_124_[10] ),
    .A1(\_122_[10] ),
    .S(_06390_),
    .X(_06393_));
 sky130_fd_sc_hd__clkbuf_1 _12704_ (.A(_06393_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _12705_ (.A0(\_124_[11] ),
    .A1(\_122_[11] ),
    .S(_06390_),
    .X(_06394_));
 sky130_fd_sc_hd__clkbuf_1 _12706_ (.A(_06394_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _12707_ (.A0(\_124_[12] ),
    .A1(\_122_[12] ),
    .S(_06390_),
    .X(_06395_));
 sky130_fd_sc_hd__clkbuf_1 _12708_ (.A(_06395_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _12709_ (.A0(\_124_[13] ),
    .A1(\_122_[13] ),
    .S(_06390_),
    .X(_06396_));
 sky130_fd_sc_hd__clkbuf_1 _12710_ (.A(_06396_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _12711_ (.A0(\_124_[14] ),
    .A1(\_122_[14] ),
    .S(_06390_),
    .X(_06397_));
 sky130_fd_sc_hd__clkbuf_1 _12712_ (.A(_06397_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _12713_ (.A0(\_124_[15] ),
    .A1(\_122_[15] ),
    .S(_06390_),
    .X(_06398_));
 sky130_fd_sc_hd__clkbuf_1 _12714_ (.A(_06398_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _12715_ (.A0(\_124_[16] ),
    .A1(\_122_[16] ),
    .S(_06390_),
    .X(_06399_));
 sky130_fd_sc_hd__clkbuf_1 _12716_ (.A(_06399_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _12717_ (.A0(\_124_[17] ),
    .A1(\_122_[17] ),
    .S(_06390_),
    .X(_06400_));
 sky130_fd_sc_hd__clkbuf_1 _12718_ (.A(_06400_),
    .X(_01124_));
 sky130_fd_sc_hd__buf_4 _12719_ (.A(_01392_),
    .X(_06401_));
 sky130_fd_sc_hd__mux2_1 _12720_ (.A0(\_124_[18] ),
    .A1(\_122_[18] ),
    .S(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__clkbuf_1 _12721_ (.A(_06402_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _12722_ (.A0(\_124_[19] ),
    .A1(\_122_[19] ),
    .S(_06401_),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_1 _12723_ (.A(_06403_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _12724_ (.A0(\_124_[20] ),
    .A1(\_122_[20] ),
    .S(_06401_),
    .X(_06404_));
 sky130_fd_sc_hd__clkbuf_1 _12725_ (.A(_06404_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _12726_ (.A0(\_124_[21] ),
    .A1(\_122_[21] ),
    .S(_06401_),
    .X(_06405_));
 sky130_fd_sc_hd__clkbuf_1 _12727_ (.A(_06405_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _12728_ (.A0(\_124_[22] ),
    .A1(\_122_[22] ),
    .S(_06401_),
    .X(_06406_));
 sky130_fd_sc_hd__clkbuf_1 _12729_ (.A(_06406_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _12730_ (.A0(\_124_[23] ),
    .A1(\_122_[23] ),
    .S(_06401_),
    .X(_06407_));
 sky130_fd_sc_hd__clkbuf_1 _12731_ (.A(_06407_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _12732_ (.A0(\_124_[24] ),
    .A1(\_122_[24] ),
    .S(_06401_),
    .X(_06408_));
 sky130_fd_sc_hd__clkbuf_1 _12733_ (.A(_06408_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _12734_ (.A0(\_124_[25] ),
    .A1(\_122_[25] ),
    .S(_06401_),
    .X(_06409_));
 sky130_fd_sc_hd__clkbuf_1 _12735_ (.A(_06409_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _12736_ (.A0(\_124_[26] ),
    .A1(\_122_[26] ),
    .S(_06401_),
    .X(_06410_));
 sky130_fd_sc_hd__clkbuf_1 _12737_ (.A(_06410_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _12738_ (.A0(\_124_[27] ),
    .A1(\_122_[27] ),
    .S(_06401_),
    .X(_06411_));
 sky130_fd_sc_hd__clkbuf_1 _12739_ (.A(_06411_),
    .X(_01134_));
 sky130_fd_sc_hd__clkbuf_4 _12740_ (.A(_01392_),
    .X(_06412_));
 sky130_fd_sc_hd__mux2_1 _12741_ (.A0(\_124_[28] ),
    .A1(\_122_[28] ),
    .S(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__clkbuf_1 _12742_ (.A(_06413_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _12743_ (.A0(\_124_[29] ),
    .A1(\_122_[29] ),
    .S(_06412_),
    .X(_06414_));
 sky130_fd_sc_hd__clkbuf_1 _12744_ (.A(_06414_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _12745_ (.A0(\_124_[30] ),
    .A1(\_122_[30] ),
    .S(_06412_),
    .X(_06415_));
 sky130_fd_sc_hd__clkbuf_1 _12746_ (.A(_06415_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _12747_ (.A0(\_124_[31] ),
    .A1(\_122_[31] ),
    .S(_06412_),
    .X(_06416_));
 sky130_fd_sc_hd__clkbuf_1 _12748_ (.A(_06416_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _12749_ (.A0(\_122_[0] ),
    .A1(\_120_[0] ),
    .S(_06412_),
    .X(_06417_));
 sky130_fd_sc_hd__clkbuf_1 _12750_ (.A(_06417_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _12751_ (.A0(\_122_[1] ),
    .A1(\_120_[1] ),
    .S(_06412_),
    .X(_06418_));
 sky130_fd_sc_hd__clkbuf_1 _12752_ (.A(_06418_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _12753_ (.A0(\_122_[2] ),
    .A1(\_120_[2] ),
    .S(_06412_),
    .X(_06419_));
 sky130_fd_sc_hd__clkbuf_1 _12754_ (.A(_06419_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _12755_ (.A0(\_122_[3] ),
    .A1(\_120_[3] ),
    .S(_06412_),
    .X(_06420_));
 sky130_fd_sc_hd__clkbuf_1 _12756_ (.A(_06420_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _12757_ (.A0(\_122_[4] ),
    .A1(\_120_[4] ),
    .S(_06412_),
    .X(_06421_));
 sky130_fd_sc_hd__clkbuf_1 _12758_ (.A(_06421_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _12759_ (.A0(\_122_[5] ),
    .A1(\_120_[5] ),
    .S(_06412_),
    .X(_06422_));
 sky130_fd_sc_hd__clkbuf_1 _12760_ (.A(_06422_),
    .X(_01144_));
 sky130_fd_sc_hd__clkbuf_8 _12761_ (.A(_01392_),
    .X(_06423_));
 sky130_fd_sc_hd__mux2_1 _12762_ (.A0(\_122_[6] ),
    .A1(\_120_[6] ),
    .S(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__clkbuf_1 _12763_ (.A(_06424_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _12764_ (.A0(\_122_[7] ),
    .A1(\_120_[7] ),
    .S(_06423_),
    .X(_06425_));
 sky130_fd_sc_hd__clkbuf_1 _12765_ (.A(_06425_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _12766_ (.A0(\_122_[8] ),
    .A1(\_120_[8] ),
    .S(_06423_),
    .X(_06426_));
 sky130_fd_sc_hd__clkbuf_1 _12767_ (.A(_06426_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _12768_ (.A0(\_122_[9] ),
    .A1(\_120_[9] ),
    .S(_06423_),
    .X(_06427_));
 sky130_fd_sc_hd__clkbuf_1 _12769_ (.A(_06427_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _12770_ (.A0(\_122_[10] ),
    .A1(\_120_[10] ),
    .S(_06423_),
    .X(_06428_));
 sky130_fd_sc_hd__clkbuf_1 _12771_ (.A(_06428_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _12772_ (.A0(\_122_[11] ),
    .A1(\_120_[11] ),
    .S(_06423_),
    .X(_06429_));
 sky130_fd_sc_hd__clkbuf_1 _12773_ (.A(_06429_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _12774_ (.A0(\_122_[12] ),
    .A1(\_120_[12] ),
    .S(_06423_),
    .X(_06430_));
 sky130_fd_sc_hd__clkbuf_1 _12775_ (.A(_06430_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _12776_ (.A0(\_122_[13] ),
    .A1(\_120_[13] ),
    .S(_06423_),
    .X(_06431_));
 sky130_fd_sc_hd__clkbuf_1 _12777_ (.A(_06431_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _12778_ (.A0(\_122_[14] ),
    .A1(\_120_[14] ),
    .S(_06423_),
    .X(_06432_));
 sky130_fd_sc_hd__clkbuf_1 _12779_ (.A(_06432_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _12780_ (.A0(\_122_[15] ),
    .A1(\_120_[15] ),
    .S(_06423_),
    .X(_06433_));
 sky130_fd_sc_hd__clkbuf_1 _12781_ (.A(_06433_),
    .X(_01154_));
 sky130_fd_sc_hd__buf_4 _12782_ (.A(_01392_),
    .X(_06434_));
 sky130_fd_sc_hd__mux2_1 _12783_ (.A0(\_122_[16] ),
    .A1(\_120_[16] ),
    .S(_06434_),
    .X(_06435_));
 sky130_fd_sc_hd__clkbuf_1 _12784_ (.A(_06435_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _12785_ (.A0(\_122_[17] ),
    .A1(\_120_[17] ),
    .S(_06434_),
    .X(_06436_));
 sky130_fd_sc_hd__clkbuf_1 _12786_ (.A(_06436_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _12787_ (.A0(\_122_[18] ),
    .A1(\_120_[18] ),
    .S(_06434_),
    .X(_06437_));
 sky130_fd_sc_hd__clkbuf_1 _12788_ (.A(_06437_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _12789_ (.A0(\_122_[19] ),
    .A1(\_120_[19] ),
    .S(_06434_),
    .X(_06438_));
 sky130_fd_sc_hd__clkbuf_1 _12790_ (.A(_06438_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _12791_ (.A0(\_122_[20] ),
    .A1(\_120_[20] ),
    .S(_06434_),
    .X(_06439_));
 sky130_fd_sc_hd__clkbuf_1 _12792_ (.A(_06439_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _12793_ (.A0(\_122_[21] ),
    .A1(\_120_[21] ),
    .S(_06434_),
    .X(_06440_));
 sky130_fd_sc_hd__clkbuf_1 _12794_ (.A(_06440_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _12795_ (.A0(\_122_[22] ),
    .A1(\_120_[22] ),
    .S(_06434_),
    .X(_06441_));
 sky130_fd_sc_hd__clkbuf_1 _12796_ (.A(_06441_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _12797_ (.A0(\_122_[23] ),
    .A1(\_120_[23] ),
    .S(_06434_),
    .X(_06442_));
 sky130_fd_sc_hd__clkbuf_1 _12798_ (.A(_06442_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _12799_ (.A0(\_122_[24] ),
    .A1(\_120_[24] ),
    .S(_06434_),
    .X(_06443_));
 sky130_fd_sc_hd__clkbuf_1 _12800_ (.A(_06443_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _12801_ (.A0(\_122_[25] ),
    .A1(\_120_[25] ),
    .S(_06434_),
    .X(_06444_));
 sky130_fd_sc_hd__clkbuf_1 _12802_ (.A(_06444_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _12803_ (.A0(\_122_[26] ),
    .A1(\_120_[26] ),
    .S(_01367_),
    .X(_06445_));
 sky130_fd_sc_hd__clkbuf_1 _12804_ (.A(_06445_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _12805_ (.A0(\_122_[27] ),
    .A1(\_120_[27] ),
    .S(_01367_),
    .X(_06446_));
 sky130_fd_sc_hd__clkbuf_1 _12806_ (.A(_06446_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _12807_ (.A0(\_122_[28] ),
    .A1(\_120_[28] ),
    .S(_01367_),
    .X(_06447_));
 sky130_fd_sc_hd__clkbuf_1 _12808_ (.A(_06447_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _12809_ (.A0(\_122_[29] ),
    .A1(\_120_[29] ),
    .S(_01367_),
    .X(_06448_));
 sky130_fd_sc_hd__clkbuf_1 _12810_ (.A(_06448_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _12811_ (.A0(\_122_[30] ),
    .A1(\_120_[30] ),
    .S(_01367_),
    .X(_06449_));
 sky130_fd_sc_hd__clkbuf_1 _12812_ (.A(_06449_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _12813_ (.A0(\_122_[31] ),
    .A1(\_120_[31] ),
    .S(_01367_),
    .X(_06450_));
 sky130_fd_sc_hd__clkbuf_1 _12814_ (.A(_06450_),
    .X(_01170_));
 sky130_fd_sc_hd__clkbuf_4 _12815_ (.A(_06004_),
    .X(_06451_));
 sky130_fd_sc_hd__mux2_1 _12816_ (.A0(\_118_[0] ),
    .A1(\_120_[0] ),
    .S(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__clkbuf_1 _12817_ (.A(_06452_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _12818_ (.A0(\_118_[1] ),
    .A1(\_120_[1] ),
    .S(_06451_),
    .X(_06453_));
 sky130_fd_sc_hd__clkbuf_1 _12819_ (.A(_06453_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _12820_ (.A0(\_118_[2] ),
    .A1(\_120_[2] ),
    .S(_06451_),
    .X(_06454_));
 sky130_fd_sc_hd__clkbuf_1 _12821_ (.A(_06454_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _12822_ (.A0(\_118_[3] ),
    .A1(\_120_[3] ),
    .S(_06451_),
    .X(_06455_));
 sky130_fd_sc_hd__clkbuf_1 _12823_ (.A(_06455_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _12824_ (.A0(\_118_[4] ),
    .A1(\_120_[4] ),
    .S(_06451_),
    .X(_06456_));
 sky130_fd_sc_hd__clkbuf_1 _12825_ (.A(_06456_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _12826_ (.A0(\_118_[5] ),
    .A1(\_120_[5] ),
    .S(_06451_),
    .X(_06457_));
 sky130_fd_sc_hd__clkbuf_1 _12827_ (.A(_06457_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _12828_ (.A0(\_118_[6] ),
    .A1(\_120_[6] ),
    .S(_06451_),
    .X(_06458_));
 sky130_fd_sc_hd__clkbuf_1 _12829_ (.A(_06458_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _12830_ (.A0(\_118_[7] ),
    .A1(\_120_[7] ),
    .S(_06451_),
    .X(_06459_));
 sky130_fd_sc_hd__clkbuf_1 _12831_ (.A(_06459_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _12832_ (.A0(\_118_[8] ),
    .A1(\_120_[8] ),
    .S(_06451_),
    .X(_06460_));
 sky130_fd_sc_hd__clkbuf_1 _12833_ (.A(_06460_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _12834_ (.A0(\_118_[9] ),
    .A1(\_120_[9] ),
    .S(_06451_),
    .X(_06461_));
 sky130_fd_sc_hd__clkbuf_1 _12835_ (.A(_06461_),
    .X(_01180_));
 sky130_fd_sc_hd__buf_4 _12836_ (.A(_06004_),
    .X(_06462_));
 sky130_fd_sc_hd__mux2_1 _12837_ (.A0(\_118_[10] ),
    .A1(\_120_[10] ),
    .S(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__clkbuf_1 _12838_ (.A(_06463_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _12839_ (.A0(\_118_[11] ),
    .A1(\_120_[11] ),
    .S(_06462_),
    .X(_06464_));
 sky130_fd_sc_hd__clkbuf_1 _12840_ (.A(_06464_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _12841_ (.A0(\_118_[12] ),
    .A1(\_120_[12] ),
    .S(_06462_),
    .X(_06465_));
 sky130_fd_sc_hd__clkbuf_1 _12842_ (.A(_06465_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _12843_ (.A0(\_118_[13] ),
    .A1(\_120_[13] ),
    .S(_06462_),
    .X(_06466_));
 sky130_fd_sc_hd__clkbuf_1 _12844_ (.A(_06466_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _12845_ (.A0(\_118_[14] ),
    .A1(\_120_[14] ),
    .S(_06462_),
    .X(_06467_));
 sky130_fd_sc_hd__clkbuf_1 _12846_ (.A(_06467_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _12847_ (.A0(\_118_[15] ),
    .A1(\_120_[15] ),
    .S(_06462_),
    .X(_06468_));
 sky130_fd_sc_hd__clkbuf_1 _12848_ (.A(_06468_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _12849_ (.A0(\_118_[16] ),
    .A1(\_120_[16] ),
    .S(_06462_),
    .X(_06469_));
 sky130_fd_sc_hd__clkbuf_1 _12850_ (.A(_06469_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _12851_ (.A0(\_118_[17] ),
    .A1(\_120_[17] ),
    .S(_06462_),
    .X(_06470_));
 sky130_fd_sc_hd__clkbuf_1 _12852_ (.A(_06470_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _12853_ (.A0(\_118_[18] ),
    .A1(\_120_[18] ),
    .S(_06462_),
    .X(_06471_));
 sky130_fd_sc_hd__clkbuf_1 _12854_ (.A(_06471_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _12855_ (.A0(\_118_[19] ),
    .A1(\_120_[19] ),
    .S(_06462_),
    .X(_06472_));
 sky130_fd_sc_hd__clkbuf_1 _12856_ (.A(_06472_),
    .X(_01190_));
 sky130_fd_sc_hd__clkbuf_4 _12857_ (.A(_06004_),
    .X(_06473_));
 sky130_fd_sc_hd__mux2_1 _12858_ (.A0(\_118_[20] ),
    .A1(\_120_[20] ),
    .S(_06473_),
    .X(_06474_));
 sky130_fd_sc_hd__clkbuf_1 _12859_ (.A(_06474_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _12860_ (.A0(\_118_[21] ),
    .A1(\_120_[21] ),
    .S(_06473_),
    .X(_06475_));
 sky130_fd_sc_hd__clkbuf_1 _12861_ (.A(_06475_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _12862_ (.A0(\_118_[22] ),
    .A1(\_120_[22] ),
    .S(_06473_),
    .X(_06476_));
 sky130_fd_sc_hd__clkbuf_1 _12863_ (.A(_06476_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _12864_ (.A0(\_118_[23] ),
    .A1(\_120_[23] ),
    .S(_06473_),
    .X(_06477_));
 sky130_fd_sc_hd__clkbuf_1 _12865_ (.A(_06477_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _12866_ (.A0(\_118_[24] ),
    .A1(\_120_[24] ),
    .S(_06473_),
    .X(_06478_));
 sky130_fd_sc_hd__clkbuf_1 _12867_ (.A(_06478_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _12868_ (.A0(\_118_[25] ),
    .A1(\_120_[25] ),
    .S(_06473_),
    .X(_06479_));
 sky130_fd_sc_hd__clkbuf_1 _12869_ (.A(_06479_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _12870_ (.A0(\_118_[26] ),
    .A1(\_120_[26] ),
    .S(_06473_),
    .X(_06480_));
 sky130_fd_sc_hd__clkbuf_1 _12871_ (.A(_06480_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _12872_ (.A0(\_118_[27] ),
    .A1(\_120_[27] ),
    .S(_06473_),
    .X(_06481_));
 sky130_fd_sc_hd__clkbuf_1 _12873_ (.A(_06481_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _12874_ (.A0(\_118_[28] ),
    .A1(\_120_[28] ),
    .S(_06473_),
    .X(_06482_));
 sky130_fd_sc_hd__clkbuf_1 _12875_ (.A(_06482_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _12876_ (.A0(\_118_[29] ),
    .A1(\_120_[29] ),
    .S(_06473_),
    .X(_06483_));
 sky130_fd_sc_hd__clkbuf_1 _12877_ (.A(_06483_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _12878_ (.A0(\_118_[30] ),
    .A1(\_120_[30] ),
    .S(_01361_),
    .X(_06484_));
 sky130_fd_sc_hd__clkbuf_1 _12879_ (.A(_06484_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _12880_ (.A0(\_118_[31] ),
    .A1(\_120_[31] ),
    .S(_01361_),
    .X(_06485_));
 sky130_fd_sc_hd__clkbuf_1 _12881_ (.A(_06485_),
    .X(_01202_));
 sky130_fd_sc_hd__or2_1 _12882_ (.A(_099_),
    .B(_05190_),
    .X(_06486_));
 sky130_fd_sc_hd__o211a_1 _12883_ (.A1(net25),
    .A2(_05196_),
    .B1(_06486_),
    .C1(_01425_),
    .X(_01203_));
 sky130_fd_sc_hd__and3_1 _12884_ (.A(_01276_),
    .B(_01292_),
    .C(_03958_),
    .X(_06487_));
 sky130_fd_sc_hd__a32o_1 _12885_ (.A1(_01233_),
    .A2(_01239_),
    .A3(_06487_),
    .B1(_01296_),
    .B2(_096_),
    .X(_06488_));
 sky130_fd_sc_hd__and2_1 _12886_ (.A(_03864_),
    .B(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__clkbuf_1 _12887_ (.A(_06489_),
    .X(_01204_));
 sky130_fd_sc_hd__a22o_1 _12888_ (.A1(_093_),
    .A2(_01296_),
    .B1(_04060_),
    .B2(_06487_),
    .X(_06490_));
 sky130_fd_sc_hd__and2_1 _12889_ (.A(_04648_),
    .B(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__clkbuf_1 _12890_ (.A(_06491_),
    .X(_01205_));
 sky130_fd_sc_hd__dfxtp_1 _12891_ (.CLK(clknet_leaf_68_clk),
    .D(_00115_),
    .Q(\_116_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12892_ (.CLK(clknet_leaf_68_clk),
    .D(_00116_),
    .Q(\_116_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12893_ (.CLK(clknet_leaf_68_clk),
    .D(_00117_),
    .Q(\_116_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12894_ (.CLK(clknet_leaf_71_clk),
    .D(_00118_),
    .Q(\_116_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12895_ (.CLK(clknet_leaf_72_clk),
    .D(_00119_),
    .Q(\_116_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12896_ (.CLK(clknet_leaf_72_clk),
    .D(_00120_),
    .Q(\_116_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12897_ (.CLK(clknet_leaf_73_clk),
    .D(_00121_),
    .Q(\_116_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12898_ (.CLK(clknet_leaf_73_clk),
    .D(_00122_),
    .Q(\_116_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12899_ (.CLK(clknet_leaf_89_clk),
    .D(_00123_),
    .Q(\_116_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12900_ (.CLK(clknet_leaf_72_clk),
    .D(_00124_),
    .Q(\_116_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12901_ (.CLK(clknet_leaf_90_clk),
    .D(_00125_),
    .Q(\_116_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12902_ (.CLK(clknet_leaf_91_clk),
    .D(_00126_),
    .Q(\_116_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12903_ (.CLK(clknet_leaf_91_clk),
    .D(_00127_),
    .Q(\_116_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12904_ (.CLK(clknet_leaf_93_clk),
    .D(_00128_),
    .Q(\_116_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12905_ (.CLK(clknet_leaf_93_clk),
    .D(_00129_),
    .Q(\_116_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12906_ (.CLK(clknet_leaf_86_clk),
    .D(_00130_),
    .Q(\_116_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12907_ (.CLK(clknet_leaf_86_clk),
    .D(_00131_),
    .Q(\_116_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12908_ (.CLK(clknet_leaf_86_clk),
    .D(_00132_),
    .Q(\_116_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12909_ (.CLK(clknet_leaf_86_clk),
    .D(_00133_),
    .Q(\_116_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12910_ (.CLK(clknet_leaf_89_clk),
    .D(_00134_),
    .Q(\_116_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12911_ (.CLK(clknet_leaf_74_clk),
    .D(_00135_),
    .Q(\_116_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12912_ (.CLK(clknet_leaf_88_clk),
    .D(_00136_),
    .Q(\_116_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12913_ (.CLK(clknet_leaf_88_clk),
    .D(_00137_),
    .Q(\_116_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12914_ (.CLK(clknet_leaf_88_clk),
    .D(_00138_),
    .Q(\_116_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12915_ (.CLK(clknet_leaf_88_clk),
    .D(_00139_),
    .Q(\_116_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12916_ (.CLK(clknet_leaf_88_clk),
    .D(_00140_),
    .Q(\_116_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12917_ (.CLK(clknet_leaf_88_clk),
    .D(_00141_),
    .Q(\_116_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12918_ (.CLK(clknet_leaf_87_clk),
    .D(_00142_),
    .Q(\_116_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12919_ (.CLK(clknet_leaf_73_clk),
    .D(_00143_),
    .Q(\_116_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12920_ (.CLK(clknet_leaf_73_clk),
    .D(_00144_),
    .Q(\_116_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12921_ (.CLK(clknet_leaf_73_clk),
    .D(_00145_),
    .Q(\_116_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12922_ (.CLK(clknet_leaf_88_clk),
    .D(_00146_),
    .Q(\_116_[31] ));
 sky130_fd_sc_hd__dfrtp_2 _12923_ (.CLK(clknet_leaf_32_clk),
    .D(\_436_[0] ),
    .RESET_B(_00100_),
    .Q(\_392_[0] ));
 sky130_fd_sc_hd__dfstp_2 _12924_ (.CLK(clknet_leaf_28_clk),
    .D(\_436_[1] ),
    .SET_B(_00101_),
    .Q(\_392_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12925_ (.CLK(clknet_leaf_32_clk),
    .D(\_436_[2] ),
    .RESET_B(_00102_),
    .Q(\_392_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12926_ (.CLK(clknet_leaf_31_clk),
    .D(\_436_[3] ),
    .RESET_B(_00103_),
    .Q(\_392_[3] ));
 sky130_fd_sc_hd__dfstp_2 _12927_ (.CLK(clknet_leaf_30_clk),
    .D(\_436_[4] ),
    .SET_B(_00104_),
    .Q(\_392_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12928_ (.CLK(clknet_leaf_40_clk),
    .D(_00147_),
    .Q(\_246_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12929_ (.CLK(clknet_leaf_41_clk),
    .D(_00148_),
    .Q(\_246_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12930_ (.CLK(clknet_leaf_41_clk),
    .D(_00149_),
    .Q(\_246_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12931_ (.CLK(clknet_leaf_40_clk),
    .D(_00150_),
    .Q(\_246_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12932_ (.CLK(clknet_leaf_39_clk),
    .D(_00151_),
    .Q(\_246_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12933_ (.CLK(clknet_leaf_39_clk),
    .D(_00152_),
    .Q(\_246_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12934_ (.CLK(clknet_leaf_39_clk),
    .D(_00153_),
    .Q(\_246_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12935_ (.CLK(clknet_leaf_40_clk),
    .D(_00154_),
    .Q(\_246_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12936_ (.CLK(clknet_leaf_40_clk),
    .D(_00155_),
    .Q(\_246_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12937_ (.CLK(clknet_leaf_39_clk),
    .D(_00156_),
    .Q(\_246_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12938_ (.CLK(clknet_leaf_21_clk),
    .D(_00157_),
    .Q(\_246_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12939_ (.CLK(clknet_leaf_21_clk),
    .D(_00158_),
    .Q(\_246_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12940_ (.CLK(clknet_leaf_40_clk),
    .D(_00159_),
    .Q(\_246_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12941_ (.CLK(clknet_leaf_39_clk),
    .D(_00160_),
    .Q(\_246_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12942_ (.CLK(clknet_leaf_39_clk),
    .D(_00161_),
    .Q(\_246_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12943_ (.CLK(clknet_leaf_21_clk),
    .D(_00162_),
    .Q(\_246_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12944_ (.CLK(clknet_leaf_39_clk),
    .D(_00163_),
    .Q(\_246_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12945_ (.CLK(clknet_leaf_21_clk),
    .D(_00164_),
    .Q(\_246_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12946_ (.CLK(clknet_leaf_21_clk),
    .D(_00165_),
    .Q(\_246_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12947_ (.CLK(clknet_leaf_30_clk),
    .D(_00166_),
    .Q(\_246_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12948_ (.CLK(clknet_leaf_30_clk),
    .D(_00167_),
    .Q(\_246_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12949_ (.CLK(clknet_leaf_29_clk),
    .D(_00168_),
    .Q(\_246_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12950_ (.CLK(clknet_leaf_29_clk),
    .D(_00169_),
    .Q(\_246_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12951_ (.CLK(clknet_leaf_22_clk),
    .D(_00170_),
    .Q(\_246_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12952_ (.CLK(clknet_leaf_21_clk),
    .D(_00171_),
    .Q(\_246_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12953_ (.CLK(clknet_leaf_21_clk),
    .D(_00172_),
    .Q(\_246_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12954_ (.CLK(clknet_leaf_30_clk),
    .D(_00173_),
    .Q(\_246_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12955_ (.CLK(clknet_leaf_21_clk),
    .D(_00174_),
    .Q(\_246_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12956_ (.CLK(clknet_leaf_21_clk),
    .D(_00175_),
    .Q(\_246_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12957_ (.CLK(clknet_leaf_21_clk),
    .D(_00176_),
    .Q(\_246_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12958_ (.CLK(clknet_leaf_22_clk),
    .D(_00177_),
    .Q(\_246_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12959_ (.CLK(clknet_leaf_20_clk),
    .D(_00178_),
    .Q(\_246_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12960_ (.CLK(clknet_leaf_43_clk),
    .D(_00179_),
    .Q(\_243_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12961_ (.CLK(clknet_leaf_20_clk),
    .D(_00180_),
    .Q(\_243_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12962_ (.CLK(clknet_leaf_39_clk),
    .D(_00181_),
    .Q(\_243_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12963_ (.CLK(clknet_leaf_40_clk),
    .D(_00182_),
    .Q(\_243_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12964_ (.CLK(clknet_leaf_20_clk),
    .D(_00183_),
    .Q(\_243_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12965_ (.CLK(clknet_leaf_19_clk),
    .D(_00184_),
    .Q(\_243_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12966_ (.CLK(clknet_leaf_20_clk),
    .D(_00185_),
    .Q(\_243_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12967_ (.CLK(clknet_leaf_17_clk),
    .D(_00186_),
    .Q(\_243_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12968_ (.CLK(clknet_leaf_43_clk),
    .D(_00187_),
    .Q(\_243_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12969_ (.CLK(clknet_leaf_20_clk),
    .D(_00188_),
    .Q(\_243_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12970_ (.CLK(clknet_leaf_19_clk),
    .D(_00189_),
    .Q(\_243_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12971_ (.CLK(clknet_leaf_18_clk),
    .D(_00190_),
    .Q(\_243_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12972_ (.CLK(clknet_leaf_17_clk),
    .D(_00191_),
    .Q(\_243_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12973_ (.CLK(clknet_leaf_19_clk),
    .D(_00192_),
    .Q(\_243_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12974_ (.CLK(clknet_leaf_18_clk),
    .D(_00193_),
    .Q(\_243_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12975_ (.CLK(clknet_leaf_18_clk),
    .D(_00194_),
    .Q(\_243_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12976_ (.CLK(clknet_leaf_14_clk),
    .D(_00195_),
    .Q(\_243_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12977_ (.CLK(clknet_leaf_14_clk),
    .D(_00196_),
    .Q(\_243_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12978_ (.CLK(clknet_leaf_23_clk),
    .D(_00197_),
    .Q(\_243_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12979_ (.CLK(clknet_leaf_23_clk),
    .D(_00198_),
    .Q(\_243_[19] ));
 sky130_fd_sc_hd__dfxtp_2 _12980_ (.CLK(clknet_leaf_23_clk),
    .D(_00199_),
    .Q(\_243_[20] ));
 sky130_fd_sc_hd__dfxtp_2 _12981_ (.CLK(clknet_leaf_23_clk),
    .D(_00200_),
    .Q(\_243_[21] ));
 sky130_fd_sc_hd__dfxtp_2 _12982_ (.CLK(clknet_leaf_23_clk),
    .D(_00201_),
    .Q(\_243_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12983_ (.CLK(clknet_leaf_10_clk),
    .D(_00202_),
    .Q(\_243_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12984_ (.CLK(clknet_leaf_14_clk),
    .D(_00203_),
    .Q(\_243_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12985_ (.CLK(clknet_leaf_14_clk),
    .D(_00204_),
    .Q(\_243_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12986_ (.CLK(clknet_leaf_13_clk),
    .D(_00205_),
    .Q(\_243_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12987_ (.CLK(clknet_leaf_13_clk),
    .D(_00206_),
    .Q(\_243_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12988_ (.CLK(clknet_leaf_13_clk),
    .D(_00207_),
    .Q(\_243_[28] ));
 sky130_fd_sc_hd__dfxtp_2 _12989_ (.CLK(clknet_leaf_22_clk),
    .D(_00208_),
    .Q(\_243_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12990_ (.CLK(clknet_leaf_22_clk),
    .D(_00209_),
    .Q(\_243_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12991_ (.CLK(clknet_leaf_19_clk),
    .D(_00210_),
    .Q(\_243_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12992_ (.CLK(clknet_leaf_17_clk),
    .D(_00211_),
    .Q(\_240_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12993_ (.CLK(clknet_leaf_17_clk),
    .D(_00212_),
    .Q(\_240_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12994_ (.CLK(clknet_leaf_15_clk),
    .D(_00213_),
    .Q(\_240_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12995_ (.CLK(clknet_leaf_15_clk),
    .D(_00214_),
    .Q(\_240_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12996_ (.CLK(clknet_leaf_20_clk),
    .D(_00215_),
    .Q(\_240_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12997_ (.CLK(clknet_leaf_19_clk),
    .D(_00216_),
    .Q(\_240_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12998_ (.CLK(clknet_leaf_22_clk),
    .D(_00217_),
    .Q(\_240_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12999_ (.CLK(clknet_leaf_15_clk),
    .D(_00218_),
    .Q(\_240_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13000_ (.CLK(clknet_leaf_19_clk),
    .D(_00219_),
    .Q(\_240_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13001_ (.CLK(clknet_leaf_20_clk),
    .D(_00220_),
    .Q(\_240_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13002_ (.CLK(clknet_leaf_19_clk),
    .D(_00221_),
    .Q(\_240_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13003_ (.CLK(clknet_leaf_14_clk),
    .D(_00222_),
    .Q(\_240_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13004_ (.CLK(clknet_leaf_17_clk),
    .D(_00223_),
    .Q(\_240_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13005_ (.CLK(clknet_leaf_14_clk),
    .D(_00224_),
    .Q(\_240_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13006_ (.CLK(clknet_leaf_14_clk),
    .D(_00225_),
    .Q(\_240_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13007_ (.CLK(clknet_leaf_18_clk),
    .D(_00226_),
    .Q(\_240_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13008_ (.CLK(clknet_leaf_14_clk),
    .D(_00227_),
    .Q(\_240_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13009_ (.CLK(clknet_leaf_10_clk),
    .D(_00228_),
    .Q(\_240_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13010_ (.CLK(clknet_leaf_14_clk),
    .D(_00229_),
    .Q(\_240_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13011_ (.CLK(clknet_leaf_9_clk),
    .D(_00230_),
    .Q(\_240_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13012_ (.CLK(clknet_leaf_3_clk),
    .D(_00231_),
    .Q(\_240_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13013_ (.CLK(clknet_leaf_3_clk),
    .D(_00232_),
    .Q(\_240_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13014_ (.CLK(clknet_leaf_3_clk),
    .D(_00233_),
    .Q(\_240_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13015_ (.CLK(clknet_leaf_3_clk),
    .D(_00234_),
    .Q(\_240_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13016_ (.CLK(clknet_leaf_14_clk),
    .D(_00235_),
    .Q(\_240_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13017_ (.CLK(clknet_leaf_14_clk),
    .D(_00236_),
    .Q(\_240_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13018_ (.CLK(clknet_leaf_12_clk),
    .D(_00237_),
    .Q(\_240_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13019_ (.CLK(clknet_leaf_13_clk),
    .D(_00238_),
    .Q(\_240_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13020_ (.CLK(clknet_leaf_13_clk),
    .D(_00239_),
    .Q(\_240_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13021_ (.CLK(clknet_leaf_3_clk),
    .D(_00240_),
    .Q(\_240_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13022_ (.CLK(clknet_leaf_11_clk),
    .D(_00241_),
    .Q(\_240_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13023_ (.CLK(clknet_leaf_13_clk),
    .D(_00242_),
    .Q(\_240_[31] ));
 sky130_fd_sc_hd__dfxtp_4 _13024_ (.CLK(clknet_leaf_17_clk),
    .D(_00243_),
    .Q(\_237_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13025_ (.CLK(clknet_leaf_17_clk),
    .D(_00244_),
    .Q(\_237_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13026_ (.CLK(clknet_leaf_17_clk),
    .D(_00245_),
    .Q(\_237_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13027_ (.CLK(clknet_leaf_17_clk),
    .D(_00246_),
    .Q(\_237_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13028_ (.CLK(clknet_leaf_43_clk),
    .D(_00247_),
    .Q(\_237_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13029_ (.CLK(clknet_leaf_42_clk),
    .D(_00248_),
    .Q(\_237_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13030_ (.CLK(clknet_leaf_42_clk),
    .D(_00249_),
    .Q(\_237_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13031_ (.CLK(clknet_leaf_43_clk),
    .D(_00250_),
    .Q(\_237_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13032_ (.CLK(clknet_leaf_42_clk),
    .D(_00251_),
    .Q(\_237_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13033_ (.CLK(clknet_leaf_42_clk),
    .D(_00252_),
    .Q(\_237_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13034_ (.CLK(clknet_leaf_45_clk),
    .D(_00253_),
    .Q(\_237_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13035_ (.CLK(clknet_leaf_45_clk),
    .D(_00254_),
    .Q(\_237_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13036_ (.CLK(clknet_opt_1_0_clk),
    .D(_00255_),
    .Q(\_237_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13037_ (.CLK(clknet_leaf_81_clk),
    .D(_00256_),
    .Q(\_237_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13038_ (.CLK(clknet_4_9_0_clk),
    .D(_00257_),
    .Q(\_237_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13039_ (.CLK(clknet_4_9_0_clk),
    .D(_00258_),
    .Q(\_237_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13040_ (.CLK(clknet_leaf_83_clk),
    .D(_00259_),
    .Q(\_237_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13041_ (.CLK(clknet_leaf_110_clk),
    .D(_00260_),
    .Q(\_237_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13042_ (.CLK(clknet_leaf_110_clk),
    .D(_00261_),
    .Q(\_237_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13043_ (.CLK(clknet_leaf_110_clk),
    .D(_00262_),
    .Q(\_237_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13044_ (.CLK(clknet_leaf_108_clk),
    .D(_00263_),
    .Q(\_237_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13045_ (.CLK(clknet_leaf_108_clk),
    .D(_00264_),
    .Q(\_237_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13046_ (.CLK(clknet_leaf_108_clk),
    .D(_00265_),
    .Q(\_237_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13047_ (.CLK(clknet_leaf_109_clk),
    .D(_00266_),
    .Q(\_237_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13048_ (.CLK(clknet_leaf_110_clk),
    .D(_00267_),
    .Q(\_237_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13049_ (.CLK(clknet_leaf_85_clk),
    .D(_00268_),
    .Q(\_237_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13050_ (.CLK(clknet_leaf_108_clk),
    .D(_00269_),
    .Q(\_237_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13051_ (.CLK(clknet_leaf_85_clk),
    .D(_00270_),
    .Q(\_237_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13052_ (.CLK(clknet_leaf_110_clk),
    .D(_00271_),
    .Q(\_237_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13053_ (.CLK(clknet_leaf_108_clk),
    .D(_00272_),
    .Q(\_237_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13054_ (.CLK(clknet_leaf_110_clk),
    .D(_00273_),
    .Q(\_237_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13055_ (.CLK(clknet_leaf_85_clk),
    .D(_00274_),
    .Q(\_237_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13056_ (.CLK(clknet_leaf_13_clk),
    .D(_00275_),
    .Q(\_234_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13057_ (.CLK(clknet_leaf_15_clk),
    .D(_00276_),
    .Q(\_234_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13058_ (.CLK(clknet_leaf_112_clk),
    .D(_00277_),
    .Q(\_234_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13059_ (.CLK(clknet_leaf_15_clk),
    .D(_00278_),
    .Q(\_234_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13060_ (.CLK(clknet_leaf_110_clk),
    .D(_00279_),
    .Q(\_234_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13061_ (.CLK(clknet_leaf_110_clk),
    .D(_00280_),
    .Q(\_234_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13062_ (.CLK(clknet_leaf_112_clk),
    .D(_00281_),
    .Q(\_234_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13063_ (.CLK(clknet_leaf_109_clk),
    .D(_00282_),
    .Q(\_234_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13064_ (.CLK(clknet_leaf_110_clk),
    .D(_00283_),
    .Q(\_234_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13065_ (.CLK(clknet_leaf_109_clk),
    .D(_00284_),
    .Q(\_234_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13066_ (.CLK(clknet_leaf_110_clk),
    .D(_00285_),
    .Q(\_234_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13067_ (.CLK(clknet_leaf_106_clk),
    .D(_00286_),
    .Q(\_234_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13068_ (.CLK(clknet_leaf_83_clk),
    .D(_00287_),
    .Q(\_234_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13069_ (.CLK(clknet_leaf_83_clk),
    .D(_00288_),
    .Q(\_234_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13070_ (.CLK(clknet_leaf_83_clk),
    .D(_00289_),
    .Q(\_234_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13071_ (.CLK(clknet_leaf_107_clk),
    .D(_00290_),
    .Q(\_234_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13072_ (.CLK(clknet_leaf_99_clk),
    .D(_00291_),
    .Q(\_234_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13073_ (.CLK(clknet_leaf_99_clk),
    .D(_00292_),
    .Q(\_234_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13074_ (.CLK(clknet_leaf_99_clk),
    .D(_00293_),
    .Q(\_234_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13075_ (.CLK(clknet_leaf_99_clk),
    .D(_00294_),
    .Q(\_234_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13076_ (.CLK(clknet_leaf_99_clk),
    .D(_00295_),
    .Q(\_234_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13077_ (.CLK(clknet_leaf_100_clk),
    .D(_00296_),
    .Q(\_234_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13078_ (.CLK(clknet_leaf_101_clk),
    .D(_00297_),
    .Q(\_234_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13079_ (.CLK(clknet_leaf_100_clk),
    .D(_00298_),
    .Q(\_234_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13080_ (.CLK(clknet_leaf_100_clk),
    .D(_00299_),
    .Q(\_234_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13081_ (.CLK(clknet_leaf_99_clk),
    .D(_00300_),
    .Q(\_234_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13082_ (.CLK(clknet_leaf_102_clk),
    .D(_00301_),
    .Q(\_234_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13083_ (.CLK(clknet_leaf_107_clk),
    .D(_00302_),
    .Q(\_234_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13084_ (.CLK(clknet_leaf_100_clk),
    .D(_00303_),
    .Q(\_234_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13085_ (.CLK(clknet_leaf_102_clk),
    .D(_00304_),
    .Q(\_234_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13086_ (.CLK(clknet_leaf_104_clk),
    .D(_00305_),
    .Q(\_234_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13087_ (.CLK(clknet_leaf_104_clk),
    .D(_00306_),
    .Q(\_234_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13088_ (.CLK(clknet_leaf_115_clk),
    .D(_00307_),
    .Q(\_231_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13089_ (.CLK(clknet_leaf_111_clk),
    .D(_00308_),
    .Q(\_231_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13090_ (.CLK(clknet_leaf_115_clk),
    .D(_00309_),
    .Q(\_231_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13091_ (.CLK(clknet_leaf_115_clk),
    .D(_00310_),
    .Q(\_231_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13092_ (.CLK(clknet_leaf_111_clk),
    .D(_00311_),
    .Q(\_231_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13093_ (.CLK(clknet_leaf_111_clk),
    .D(_00312_),
    .Q(\_231_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13094_ (.CLK(clknet_leaf_111_clk),
    .D(_00313_),
    .Q(\_231_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13095_ (.CLK(clknet_leaf_106_clk),
    .D(_00314_),
    .Q(\_231_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13096_ (.CLK(clknet_leaf_109_clk),
    .D(_00315_),
    .Q(\_231_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13097_ (.CLK(clknet_leaf_116_clk),
    .D(_00316_),
    .Q(\_231_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13098_ (.CLK(clknet_leaf_106_clk),
    .D(_00317_),
    .Q(\_231_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13099_ (.CLK(clknet_leaf_106_clk),
    .D(_00318_),
    .Q(\_231_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13100_ (.CLK(clknet_leaf_109_clk),
    .D(_00319_),
    .Q(\_231_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13101_ (.CLK(clknet_leaf_116_clk),
    .D(_00320_),
    .Q(\_231_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13102_ (.CLK(clknet_leaf_116_clk),
    .D(_00321_),
    .Q(\_231_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13103_ (.CLK(clknet_leaf_117_clk),
    .D(_00322_),
    .Q(\_231_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13104_ (.CLK(clknet_leaf_105_clk),
    .D(_00323_),
    .Q(\_231_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13105_ (.CLK(clknet_leaf_117_clk),
    .D(_00324_),
    .Q(\_231_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13106_ (.CLK(clknet_leaf_117_clk),
    .D(_00325_),
    .Q(\_231_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13107_ (.CLK(clknet_leaf_118_clk),
    .D(_00326_),
    .Q(\_231_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13108_ (.CLK(clknet_leaf_104_clk),
    .D(_00327_),
    .Q(\_231_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13109_ (.CLK(clknet_leaf_118_clk),
    .D(_00328_),
    .Q(\_231_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13110_ (.CLK(clknet_leaf_118_clk),
    .D(_00329_),
    .Q(\_231_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13111_ (.CLK(clknet_leaf_103_clk),
    .D(_00330_),
    .Q(\_231_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13112_ (.CLK(clknet_leaf_103_clk),
    .D(_00331_),
    .Q(\_231_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13113_ (.CLK(clknet_leaf_103_clk),
    .D(_00332_),
    .Q(\_231_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13114_ (.CLK(clknet_leaf_119_clk),
    .D(_00333_),
    .Q(\_231_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13115_ (.CLK(clknet_leaf_120_clk),
    .D(_00334_),
    .Q(\_231_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13116_ (.CLK(clknet_leaf_119_clk),
    .D(_00335_),
    .Q(\_231_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13117_ (.CLK(clknet_leaf_119_clk),
    .D(_00336_),
    .Q(\_231_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13118_ (.CLK(clknet_leaf_103_clk),
    .D(_00337_),
    .Q(\_231_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13119_ (.CLK(clknet_leaf_119_clk),
    .D(_00338_),
    .Q(\_231_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13120_ (.CLK(clknet_leaf_117_clk),
    .D(_00339_),
    .Q(\_228_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13121_ (.CLK(clknet_leaf_112_clk),
    .D(_00340_),
    .Q(\_228_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13122_ (.CLK(clknet_leaf_115_clk),
    .D(_00341_),
    .Q(\_228_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13123_ (.CLK(clknet_leaf_116_clk),
    .D(_00342_),
    .Q(\_228_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13124_ (.CLK(clknet_leaf_112_clk),
    .D(_00343_),
    .Q(\_228_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13125_ (.CLK(clknet_leaf_111_clk),
    .D(_00344_),
    .Q(\_228_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13126_ (.CLK(clknet_leaf_109_clk),
    .D(_00345_),
    .Q(\_228_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13127_ (.CLK(clknet_leaf_106_clk),
    .D(_00346_),
    .Q(\_228_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13128_ (.CLK(clknet_leaf_111_clk),
    .D(_00347_),
    .Q(\_228_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13129_ (.CLK(clknet_leaf_117_clk),
    .D(_00348_),
    .Q(\_228_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13130_ (.CLK(clknet_leaf_106_clk),
    .D(_00349_),
    .Q(\_228_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13131_ (.CLK(clknet_leaf_117_clk),
    .D(_00350_),
    .Q(\_228_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13132_ (.CLK(clknet_leaf_109_clk),
    .D(_00351_),
    .Q(\_228_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13133_ (.CLK(clknet_leaf_117_clk),
    .D(_00352_),
    .Q(\_228_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13134_ (.CLK(clknet_leaf_115_clk),
    .D(_00353_),
    .Q(\_228_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13135_ (.CLK(clknet_leaf_117_clk),
    .D(_00354_),
    .Q(\_228_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13136_ (.CLK(clknet_leaf_117_clk),
    .D(_00355_),
    .Q(\_228_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13137_ (.CLK(clknet_leaf_118_clk),
    .D(_00356_),
    .Q(\_228_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13138_ (.CLK(clknet_leaf_118_clk),
    .D(_00357_),
    .Q(\_228_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13139_ (.CLK(clknet_leaf_118_clk),
    .D(_00358_),
    .Q(\_228_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13140_ (.CLK(clknet_4_2_0_clk),
    .D(_00359_),
    .Q(\_228_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13141_ (.CLK(clknet_leaf_118_clk),
    .D(_00360_),
    .Q(\_228_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13142_ (.CLK(clknet_leaf_120_clk),
    .D(_00361_),
    .Q(\_228_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13143_ (.CLK(clknet_leaf_119_clk),
    .D(_00362_),
    .Q(\_228_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13144_ (.CLK(clknet_leaf_103_clk),
    .D(_00363_),
    .Q(\_228_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13145_ (.CLK(clknet_leaf_119_clk),
    .D(_00364_),
    .Q(\_228_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13146_ (.CLK(clknet_leaf_120_clk),
    .D(_00365_),
    .Q(\_228_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13147_ (.CLK(clknet_leaf_120_clk),
    .D(_00366_),
    .Q(\_228_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13148_ (.CLK(clknet_leaf_119_clk),
    .D(_00367_),
    .Q(\_228_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13149_ (.CLK(clknet_leaf_119_clk),
    .D(_00368_),
    .Q(\_228_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13150_ (.CLK(clknet_leaf_120_clk),
    .D(_00369_),
    .Q(\_228_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13151_ (.CLK(clknet_leaf_104_clk),
    .D(_00370_),
    .Q(\_228_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13152_ (.CLK(clknet_leaf_116_clk),
    .D(_00371_),
    .Q(\_225_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13153_ (.CLK(clknet_leaf_13_clk),
    .D(_00372_),
    .Q(\_225_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13154_ (.CLK(clknet_leaf_2_clk),
    .D(_00373_),
    .Q(\_225_[2] ));
 sky130_fd_sc_hd__dfxtp_4 _13155_ (.CLK(clknet_leaf_112_clk),
    .D(_00374_),
    .Q(\_225_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13156_ (.CLK(clknet_leaf_111_clk),
    .D(_00375_),
    .Q(\_225_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13157_ (.CLK(clknet_leaf_111_clk),
    .D(_00376_),
    .Q(\_225_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13158_ (.CLK(clknet_leaf_109_clk),
    .D(_00377_),
    .Q(\_225_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13159_ (.CLK(clknet_leaf_111_clk),
    .D(_00378_),
    .Q(\_225_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13160_ (.CLK(clknet_leaf_109_clk),
    .D(_00379_),
    .Q(\_225_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13161_ (.CLK(clknet_leaf_109_clk),
    .D(_00380_),
    .Q(\_225_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13162_ (.CLK(clknet_leaf_106_clk),
    .D(_00381_),
    .Q(\_225_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13163_ (.CLK(clknet_leaf_106_clk),
    .D(_00382_),
    .Q(\_225_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13164_ (.CLK(clknet_leaf_109_clk),
    .D(_00383_),
    .Q(\_225_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13165_ (.CLK(clknet_leaf_109_clk),
    .D(_00384_),
    .Q(\_225_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13166_ (.CLK(clknet_leaf_106_clk),
    .D(_00385_),
    .Q(\_225_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13167_ (.CLK(clknet_leaf_108_clk),
    .D(_00386_),
    .Q(\_225_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13168_ (.CLK(clknet_leaf_105_clk),
    .D(_00387_),
    .Q(\_225_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13169_ (.CLK(clknet_leaf_105_clk),
    .D(_00388_),
    .Q(\_225_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13170_ (.CLK(clknet_leaf_100_clk),
    .D(_00389_),
    .Q(\_225_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13171_ (.CLK(clknet_leaf_105_clk),
    .D(_00390_),
    .Q(\_225_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13172_ (.CLK(clknet_leaf_104_clk),
    .D(_00391_),
    .Q(\_225_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13173_ (.CLK(clknet_leaf_103_clk),
    .D(_00392_),
    .Q(\_225_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13174_ (.CLK(clknet_leaf_103_clk),
    .D(_00393_),
    .Q(\_225_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13175_ (.CLK(clknet_leaf_101_clk),
    .D(_00394_),
    .Q(\_225_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13176_ (.CLK(clknet_leaf_103_clk),
    .D(_00395_),
    .Q(\_225_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13177_ (.CLK(clknet_leaf_103_clk),
    .D(_00396_),
    .Q(\_225_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13178_ (.CLK(clknet_leaf_101_clk),
    .D(_00397_),
    .Q(\_225_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13179_ (.CLK(clknet_leaf_102_clk),
    .D(_00398_),
    .Q(\_225_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13180_ (.CLK(clknet_leaf_102_clk),
    .D(_00399_),
    .Q(\_225_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13181_ (.CLK(clknet_leaf_102_clk),
    .D(_00400_),
    .Q(\_225_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13182_ (.CLK(clknet_leaf_103_clk),
    .D(_00401_),
    .Q(\_225_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13183_ (.CLK(clknet_leaf_120_clk),
    .D(_00402_),
    .Q(\_225_[31] ));
 sky130_fd_sc_hd__dfrtp_2 _13184_ (.CLK(clknet_leaf_31_clk),
    .D(_00403_),
    .RESET_B(_00105_),
    .Q(\_195_[0] ));
 sky130_fd_sc_hd__dfrtp_2 _13185_ (.CLK(clknet_leaf_33_clk),
    .D(_00404_),
    .RESET_B(_00106_),
    .Q(\_195_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13186_ (.CLK(clknet_leaf_33_clk),
    .D(_00405_),
    .RESET_B(_00107_),
    .Q(\_195_[2] ));
 sky130_fd_sc_hd__dfrtp_4 _13187_ (.CLK(clknet_leaf_33_clk),
    .D(_00406_),
    .RESET_B(_00108_),
    .Q(\_195_[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13188_ (.CLK(clknet_leaf_33_clk),
    .D(_00407_),
    .RESET_B(_00109_),
    .Q(\_195_[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13189_ (.CLK(clknet_leaf_33_clk),
    .D(_00408_),
    .RESET_B(_00110_),
    .Q(\_195_[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13190_ (.CLK(clknet_leaf_35_clk),
    .D(_00409_),
    .Q(\_185_[0] ));
 sky130_fd_sc_hd__dfxtp_2 _13191_ (.CLK(clknet_leaf_34_clk),
    .D(_00410_),
    .Q(\_185_[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13192_ (.CLK(clknet_leaf_34_clk),
    .D(_00411_),
    .Q(\_185_[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13193_ (.CLK(clknet_leaf_34_clk),
    .D(_00412_),
    .Q(\_185_[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13194_ (.CLK(clknet_leaf_34_clk),
    .D(_00413_),
    .Q(\_185_[4] ));
 sky130_fd_sc_hd__dfxtp_4 _13195_ (.CLK(clknet_leaf_34_clk),
    .D(_00414_),
    .Q(\_185_[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13196_ (.CLK(clknet_leaf_34_clk),
    .D(_00415_),
    .Q(\_185_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13197_ (.CLK(clknet_leaf_34_clk),
    .D(_00416_),
    .Q(\_185_[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13198_ (.CLK(clknet_leaf_34_clk),
    .D(_00417_),
    .Q(\_185_[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13199_ (.CLK(clknet_leaf_34_clk),
    .D(_00418_),
    .Q(\_185_[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13200_ (.CLK(clknet_leaf_35_clk),
    .D(_00419_),
    .Q(\_185_[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13201_ (.CLK(clknet_leaf_35_clk),
    .D(_00420_),
    .Q(\_185_[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13202_ (.CLK(clknet_leaf_35_clk),
    .D(_00421_),
    .Q(\_185_[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13203_ (.CLK(clknet_leaf_36_clk),
    .D(_00422_),
    .Q(\_185_[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13204_ (.CLK(clknet_leaf_36_clk),
    .D(_00423_),
    .Q(\_185_[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13205_ (.CLK(clknet_leaf_40_clk),
    .D(_00424_),
    .Q(\_185_[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13206_ (.CLK(clknet_leaf_41_clk),
    .D(_00425_),
    .Q(\_185_[16] ));
 sky130_fd_sc_hd__dfxtp_4 _13207_ (.CLK(clknet_leaf_42_clk),
    .D(_00426_),
    .Q(\_185_[17] ));
 sky130_fd_sc_hd__dfxtp_4 _13208_ (.CLK(clknet_leaf_41_clk),
    .D(_00427_),
    .Q(\_185_[18] ));
 sky130_fd_sc_hd__dfxtp_4 _13209_ (.CLK(clknet_leaf_42_clk),
    .D(_00428_),
    .Q(\_185_[19] ));
 sky130_fd_sc_hd__dfxtp_4 _13210_ (.CLK(clknet_leaf_41_clk),
    .D(_00429_),
    .Q(\_185_[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13211_ (.CLK(clknet_leaf_41_clk),
    .D(_00430_),
    .Q(\_185_[21] ));
 sky130_fd_sc_hd__dfxtp_4 _13212_ (.CLK(clknet_leaf_37_clk),
    .D(_00431_),
    .Q(\_185_[22] ));
 sky130_fd_sc_hd__dfxtp_4 _13213_ (.CLK(clknet_leaf_41_clk),
    .D(_00432_),
    .Q(\_185_[23] ));
 sky130_fd_sc_hd__dfxtp_4 _13214_ (.CLK(clknet_leaf_37_clk),
    .D(_00433_),
    .Q(\_185_[24] ));
 sky130_fd_sc_hd__dfxtp_4 _13215_ (.CLK(clknet_leaf_37_clk),
    .D(_00434_),
    .Q(\_185_[25] ));
 sky130_fd_sc_hd__dfxtp_4 _13216_ (.CLK(clknet_leaf_37_clk),
    .D(_00435_),
    .Q(\_185_[26] ));
 sky130_fd_sc_hd__dfxtp_4 _13217_ (.CLK(clknet_leaf_38_clk),
    .D(_00436_),
    .Q(\_185_[27] ));
 sky130_fd_sc_hd__dfxtp_4 _13218_ (.CLK(clknet_leaf_38_clk),
    .D(_00437_),
    .Q(\_185_[28] ));
 sky130_fd_sc_hd__dfxtp_2 _13219_ (.CLK(clknet_leaf_41_clk),
    .D(_00438_),
    .Q(\_185_[29] ));
 sky130_fd_sc_hd__dfxtp_2 _13220_ (.CLK(clknet_leaf_37_clk),
    .D(_00439_),
    .Q(\_185_[30] ));
 sky130_fd_sc_hd__dfxtp_2 _13221_ (.CLK(clknet_leaf_38_clk),
    .D(_00440_),
    .Q(\_185_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13222_ (.CLK(clknet_leaf_24_clk),
    .D(_00441_),
    .Q(\_182_[0] ));
 sky130_fd_sc_hd__dfxtp_2 _13223_ (.CLK(clknet_leaf_28_clk),
    .D(_00442_),
    .Q(\_182_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13224_ (.CLK(clknet_leaf_28_clk),
    .D(_00443_),
    .Q(\_182_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13225_ (.CLK(clknet_leaf_24_clk),
    .D(_00444_),
    .Q(\_182_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13226_ (.CLK(clknet_leaf_27_clk),
    .D(_00445_),
    .Q(\_182_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13227_ (.CLK(clknet_leaf_29_clk),
    .D(_00446_),
    .Q(\_182_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13228_ (.CLK(clknet_leaf_28_clk),
    .D(_00447_),
    .Q(\_182_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13229_ (.CLK(clknet_leaf_29_clk),
    .D(_00448_),
    .Q(\_182_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13230_ (.CLK(clknet_leaf_27_clk),
    .D(_00449_),
    .Q(\_182_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13231_ (.CLK(clknet_leaf_27_clk),
    .D(_00450_),
    .Q(\_182_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13232_ (.CLK(clknet_leaf_27_clk),
    .D(_00451_),
    .Q(\_182_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13233_ (.CLK(clknet_leaf_25_clk),
    .D(_00452_),
    .Q(\_182_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13234_ (.CLK(clknet_leaf_26_clk),
    .D(_00453_),
    .Q(\_182_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13235_ (.CLK(clknet_leaf_25_clk),
    .D(_00454_),
    .Q(\_182_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13236_ (.CLK(clknet_leaf_7_clk),
    .D(_00455_),
    .Q(\_182_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13237_ (.CLK(clknet_leaf_25_clk),
    .D(_00456_),
    .Q(\_182_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13238_ (.CLK(clknet_leaf_25_clk),
    .D(_00457_),
    .Q(\_182_[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13239_ (.CLK(clknet_leaf_25_clk),
    .D(_00458_),
    .Q(\_182_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13240_ (.CLK(clknet_leaf_25_clk),
    .D(_00459_),
    .Q(\_182_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13241_ (.CLK(clknet_leaf_6_clk),
    .D(_00460_),
    .Q(\_182_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13242_ (.CLK(clknet_leaf_6_clk),
    .D(_00461_),
    .Q(\_182_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13243_ (.CLK(clknet_leaf_6_clk),
    .D(_00462_),
    .Q(\_182_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13244_ (.CLK(clknet_leaf_6_clk),
    .D(_00463_),
    .Q(\_182_[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13245_ (.CLK(clknet_leaf_5_clk),
    .D(_00464_),
    .Q(\_182_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13246_ (.CLK(clknet_leaf_7_clk),
    .D(_00465_),
    .Q(\_182_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13247_ (.CLK(clknet_leaf_5_clk),
    .D(_00466_),
    .Q(\_182_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13248_ (.CLK(clknet_leaf_5_clk),
    .D(_00467_),
    .Q(\_182_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13249_ (.CLK(clknet_leaf_7_clk),
    .D(_00468_),
    .Q(\_182_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13250_ (.CLK(clknet_leaf_8_clk),
    .D(_00469_),
    .Q(\_182_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13251_ (.CLK(clknet_leaf_5_clk),
    .D(_00470_),
    .Q(\_182_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13252_ (.CLK(clknet_leaf_5_clk),
    .D(_00471_),
    .Q(\_182_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13253_ (.CLK(clknet_leaf_5_clk),
    .D(_00472_),
    .Q(\_182_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13254_ (.CLK(clknet_leaf_24_clk),
    .D(_00473_),
    .Q(\_179_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13255_ (.CLK(clknet_leaf_24_clk),
    .D(_00474_),
    .Q(\_179_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13256_ (.CLK(clknet_leaf_28_clk),
    .D(_00475_),
    .Q(\_179_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13257_ (.CLK(clknet_leaf_24_clk),
    .D(_00476_),
    .Q(\_179_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13258_ (.CLK(clknet_leaf_29_clk),
    .D(_00477_),
    .Q(\_179_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13259_ (.CLK(clknet_leaf_29_clk),
    .D(_00478_),
    .Q(\_179_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13260_ (.CLK(clknet_leaf_28_clk),
    .D(_00479_),
    .Q(\_179_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13261_ (.CLK(clknet_leaf_29_clk),
    .D(_00480_),
    .Q(\_179_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13262_ (.CLK(clknet_leaf_26_clk),
    .D(_00481_),
    .Q(\_179_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13263_ (.CLK(clknet_leaf_27_clk),
    .D(_00482_),
    .Q(\_179_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13264_ (.CLK(clknet_leaf_27_clk),
    .D(_00483_),
    .Q(\_179_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13265_ (.CLK(clknet_leaf_25_clk),
    .D(_00484_),
    .Q(\_179_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13266_ (.CLK(clknet_leaf_26_clk),
    .D(_00485_),
    .Q(\_179_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13267_ (.CLK(clknet_leaf_26_clk),
    .D(_00486_),
    .Q(\_179_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13268_ (.CLK(clknet_leaf_24_clk),
    .D(_00487_),
    .Q(\_179_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13269_ (.CLK(clknet_leaf_25_clk),
    .D(_00488_),
    .Q(\_179_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13270_ (.CLK(clknet_leaf_7_clk),
    .D(_00489_),
    .Q(\_179_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13271_ (.CLK(clknet_leaf_7_clk),
    .D(_00490_),
    .Q(\_179_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13272_ (.CLK(clknet_leaf_25_clk),
    .D(_00491_),
    .Q(\_179_[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13273_ (.CLK(clknet_leaf_25_clk),
    .D(_00492_),
    .Q(\_179_[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13274_ (.CLK(clknet_leaf_4_clk),
    .D(_00493_),
    .Q(\_179_[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13275_ (.CLK(clknet_leaf_4_clk),
    .D(_00494_),
    .Q(\_179_[21] ));
 sky130_fd_sc_hd__dfxtp_2 _13276_ (.CLK(clknet_leaf_4_clk),
    .D(_00495_),
    .Q(\_179_[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13277_ (.CLK(clknet_leaf_7_clk),
    .D(_00496_),
    .Q(\_179_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13278_ (.CLK(clknet_leaf_7_clk),
    .D(_00497_),
    .Q(\_179_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13279_ (.CLK(clknet_leaf_7_clk),
    .D(_00498_),
    .Q(\_179_[25] ));
 sky130_fd_sc_hd__dfxtp_2 _13280_ (.CLK(clknet_leaf_5_clk),
    .D(_00499_),
    .Q(\_179_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13281_ (.CLK(clknet_leaf_7_clk),
    .D(_00500_),
    .Q(\_179_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13282_ (.CLK(clknet_leaf_8_clk),
    .D(_00501_),
    .Q(\_179_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13283_ (.CLK(clknet_leaf_3_clk),
    .D(_00502_),
    .Q(\_179_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13284_ (.CLK(clknet_leaf_5_clk),
    .D(_00503_),
    .Q(\_179_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13285_ (.CLK(clknet_leaf_5_clk),
    .D(_00504_),
    .Q(\_179_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13286_ (.CLK(clknet_leaf_24_clk),
    .D(_00505_),
    .Q(\_176_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13287_ (.CLK(clknet_leaf_24_clk),
    .D(_00506_),
    .Q(\_176_[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13288_ (.CLK(clknet_leaf_24_clk),
    .D(_00507_),
    .Q(\_176_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13289_ (.CLK(clknet_leaf_24_clk),
    .D(_00508_),
    .Q(\_176_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13290_ (.CLK(clknet_leaf_24_clk),
    .D(_00509_),
    .Q(\_176_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13291_ (.CLK(clknet_leaf_26_clk),
    .D(_00510_),
    .Q(\_176_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13292_ (.CLK(clknet_leaf_26_clk),
    .D(_00511_),
    .Q(\_176_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13293_ (.CLK(clknet_leaf_24_clk),
    .D(_00512_),
    .Q(\_176_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13294_ (.CLK(clknet_leaf_26_clk),
    .D(_00513_),
    .Q(\_176_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13295_ (.CLK(clknet_leaf_26_clk),
    .D(_00514_),
    .Q(\_176_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13296_ (.CLK(clknet_leaf_26_clk),
    .D(_00515_),
    .Q(\_176_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13297_ (.CLK(clknet_leaf_24_clk),
    .D(_00516_),
    .Q(\_176_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13298_ (.CLK(clknet_leaf_26_clk),
    .D(_00517_),
    .Q(\_176_[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13299_ (.CLK(clknet_leaf_23_clk),
    .D(_00518_),
    .Q(\_176_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13300_ (.CLK(clknet_leaf_9_clk),
    .D(_00519_),
    .Q(\_176_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13301_ (.CLK(clknet_leaf_25_clk),
    .D(_00520_),
    .Q(\_176_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13302_ (.CLK(clknet_leaf_8_clk),
    .D(_00521_),
    .Q(\_176_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13303_ (.CLK(clknet_leaf_7_clk),
    .D(_00522_),
    .Q(\_176_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13304_ (.CLK(clknet_leaf_9_clk),
    .D(_00523_),
    .Q(\_176_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13305_ (.CLK(clknet_leaf_6_clk),
    .D(_00524_),
    .Q(\_176_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13306_ (.CLK(clknet_leaf_4_clk),
    .D(_00525_),
    .Q(\_176_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13307_ (.CLK(clknet_leaf_4_clk),
    .D(_00526_),
    .Q(\_176_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13308_ (.CLK(clknet_leaf_4_clk),
    .D(_00527_),
    .Q(\_176_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13309_ (.CLK(clknet_leaf_4_clk),
    .D(_00528_),
    .Q(\_176_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13310_ (.CLK(clknet_leaf_8_clk),
    .D(_00529_),
    .Q(\_176_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13311_ (.CLK(clknet_leaf_8_clk),
    .D(_00530_),
    .Q(\_176_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13312_ (.CLK(clknet_leaf_5_clk),
    .D(_00531_),
    .Q(\_176_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13313_ (.CLK(clknet_leaf_8_clk),
    .D(_00532_),
    .Q(\_176_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13314_ (.CLK(clknet_leaf_10_clk),
    .D(_00533_),
    .Q(\_176_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13315_ (.CLK(clknet_leaf_4_clk),
    .D(_00534_),
    .Q(\_176_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13316_ (.CLK(clknet_leaf_5_clk),
    .D(_00535_),
    .Q(\_176_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13317_ (.CLK(clknet_leaf_10_clk),
    .D(_00536_),
    .Q(\_176_[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13318_ (.CLK(clknet_leaf_23_clk),
    .D(_00537_),
    .Q(\_173_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13319_ (.CLK(clknet_leaf_18_clk),
    .D(_00538_),
    .Q(\_173_[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13320_ (.CLK(clknet_leaf_18_clk),
    .D(_00539_),
    .Q(\_173_[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13321_ (.CLK(clknet_leaf_18_clk),
    .D(_00540_),
    .Q(\_173_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13322_ (.CLK(clknet_leaf_22_clk),
    .D(_00541_),
    .Q(\_173_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13323_ (.CLK(clknet_leaf_23_clk),
    .D(_00542_),
    .Q(\_173_[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13324_ (.CLK(clknet_leaf_22_clk),
    .D(_00543_),
    .Q(\_173_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13325_ (.CLK(clknet_leaf_22_clk),
    .D(_00544_),
    .Q(\_173_[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13326_ (.CLK(clknet_leaf_25_clk),
    .D(_00545_),
    .Q(\_173_[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13327_ (.CLK(clknet_leaf_22_clk),
    .D(_00546_),
    .Q(\_173_[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13328_ (.CLK(clknet_leaf_25_clk),
    .D(_00547_),
    .Q(\_173_[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13329_ (.CLK(clknet_leaf_25_clk),
    .D(_00548_),
    .Q(\_173_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13330_ (.CLK(clknet_leaf_23_clk),
    .D(_00549_),
    .Q(\_173_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13331_ (.CLK(clknet_leaf_23_clk),
    .D(_00550_),
    .Q(\_173_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13332_ (.CLK(clknet_leaf_9_clk),
    .D(_00551_),
    .Q(\_173_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13333_ (.CLK(clknet_leaf_23_clk),
    .D(_00552_),
    .Q(\_173_[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13334_ (.CLK(clknet_leaf_5_clk),
    .D(_00553_),
    .Q(\_173_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13335_ (.CLK(clknet_leaf_8_clk),
    .D(_00554_),
    .Q(\_173_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13336_ (.CLK(clknet_leaf_9_clk),
    .D(_00555_),
    .Q(\_173_[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13337_ (.CLK(clknet_leaf_10_clk),
    .D(_00556_),
    .Q(\_173_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13338_ (.CLK(clknet_leaf_0_clk),
    .D(_00557_),
    .Q(\_173_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13339_ (.CLK(clknet_leaf_0_clk),
    .D(_00558_),
    .Q(\_173_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13340_ (.CLK(clknet_leaf_4_clk),
    .D(_00559_),
    .Q(\_173_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13341_ (.CLK(clknet_leaf_4_clk),
    .D(_00560_),
    .Q(\_173_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13342_ (.CLK(clknet_leaf_10_clk),
    .D(_00561_),
    .Q(\_173_[24] ));
 sky130_fd_sc_hd__dfxtp_2 _13343_ (.CLK(clknet_leaf_11_clk),
    .D(_00562_),
    .Q(\_173_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13344_ (.CLK(clknet_leaf_12_clk),
    .D(_00563_),
    .Q(\_173_[26] ));
 sky130_fd_sc_hd__dfxtp_2 _13345_ (.CLK(clknet_leaf_10_clk),
    .D(_00564_),
    .Q(\_173_[27] ));
 sky130_fd_sc_hd__dfxtp_2 _13346_ (.CLK(clknet_leaf_11_clk),
    .D(_00565_),
    .Q(\_173_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13347_ (.CLK(clknet_leaf_4_clk),
    .D(_00566_),
    .Q(\_173_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13348_ (.CLK(clknet_leaf_11_clk),
    .D(_00567_),
    .Q(\_173_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13349_ (.CLK(clknet_leaf_8_clk),
    .D(_00568_),
    .Q(\_173_[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13350_ (.CLK(clknet_leaf_0_clk),
    .D(_00569_),
    .Q(\_170_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13351_ (.CLK(clknet_leaf_2_clk),
    .D(_00570_),
    .Q(\_170_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13352_ (.CLK(clknet_leaf_0_clk),
    .D(_00571_),
    .Q(\_170_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13353_ (.CLK(clknet_leaf_2_clk),
    .D(_00572_),
    .Q(\_170_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13354_ (.CLK(clknet_leaf_11_clk),
    .D(_00573_),
    .Q(\_170_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13355_ (.CLK(clknet_leaf_12_clk),
    .D(_00574_),
    .Q(\_170_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13356_ (.CLK(clknet_leaf_3_clk),
    .D(_00575_),
    .Q(\_170_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13357_ (.CLK(clknet_leaf_0_clk),
    .D(_00576_),
    .Q(\_170_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13358_ (.CLK(clknet_leaf_11_clk),
    .D(_00577_),
    .Q(\_170_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13359_ (.CLK(clknet_leaf_0_clk),
    .D(_00578_),
    .Q(\_170_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13360_ (.CLK(clknet_leaf_2_clk),
    .D(_00579_),
    .Q(\_170_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13361_ (.CLK(clknet_leaf_0_clk),
    .D(_00580_),
    .Q(\_170_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13362_ (.CLK(clknet_leaf_2_clk),
    .D(_00581_),
    .Q(\_170_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13363_ (.CLK(clknet_leaf_124_clk),
    .D(_00582_),
    .Q(\_170_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13364_ (.CLK(clknet_leaf_124_clk),
    .D(_00583_),
    .Q(\_170_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13365_ (.CLK(clknet_leaf_124_clk),
    .D(_00584_),
    .Q(\_170_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13366_ (.CLK(clknet_leaf_125_clk),
    .D(_00585_),
    .Q(\_170_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13367_ (.CLK(clknet_leaf_125_clk),
    .D(_00586_),
    .Q(\_170_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13368_ (.CLK(clknet_leaf_125_clk),
    .D(_00587_),
    .Q(\_170_[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13369_ (.CLK(clknet_leaf_125_clk),
    .D(_00588_),
    .Q(\_170_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13370_ (.CLK(clknet_leaf_130_clk),
    .D(_00589_),
    .Q(\_170_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13371_ (.CLK(clknet_leaf_130_clk),
    .D(_00590_),
    .Q(\_170_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13372_ (.CLK(clknet_leaf_126_clk),
    .D(_00591_),
    .Q(\_170_[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13373_ (.CLK(clknet_leaf_129_clk),
    .D(_00592_),
    .Q(\_170_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13374_ (.CLK(clknet_leaf_126_clk),
    .D(_00593_),
    .Q(\_170_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13375_ (.CLK(clknet_leaf_127_clk),
    .D(_00594_),
    .Q(\_170_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13376_ (.CLK(clknet_leaf_125_clk),
    .D(_00595_),
    .Q(\_170_[26] ));
 sky130_fd_sc_hd__dfxtp_2 _13377_ (.CLK(clknet_leaf_127_clk),
    .D(_00596_),
    .Q(\_170_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13378_ (.CLK(clknet_leaf_127_clk),
    .D(_00597_),
    .Q(\_170_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13379_ (.CLK(clknet_leaf_126_clk),
    .D(_00598_),
    .Q(\_170_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13380_ (.CLK(clknet_leaf_128_clk),
    .D(_00599_),
    .Q(\_170_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13381_ (.CLK(clknet_leaf_125_clk),
    .D(_00600_),
    .Q(\_170_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13382_ (.CLK(clknet_leaf_0_clk),
    .D(_00601_),
    .Q(\_167_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13383_ (.CLK(clknet_leaf_12_clk),
    .D(_00602_),
    .Q(\_167_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13384_ (.CLK(clknet_leaf_1_clk),
    .D(_00603_),
    .Q(\_167_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13385_ (.CLK(clknet_leaf_1_clk),
    .D(_00604_),
    .Q(\_167_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13386_ (.CLK(clknet_leaf_11_clk),
    .D(_00605_),
    .Q(\_167_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13387_ (.CLK(clknet_leaf_12_clk),
    .D(_00606_),
    .Q(\_167_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13388_ (.CLK(clknet_leaf_12_clk),
    .D(_00607_),
    .Q(\_167_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13389_ (.CLK(clknet_leaf_1_clk),
    .D(_00608_),
    .Q(\_167_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13390_ (.CLK(clknet_leaf_12_clk),
    .D(_00609_),
    .Q(\_167_[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13391_ (.CLK(clknet_leaf_2_clk),
    .D(_00610_),
    .Q(\_167_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13392_ (.CLK(clknet_leaf_1_clk),
    .D(_00611_),
    .Q(\_167_[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13393_ (.CLK(clknet_leaf_130_clk),
    .D(_00612_),
    .Q(\_167_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13394_ (.CLK(clknet_leaf_124_clk),
    .D(_00613_),
    .Q(\_167_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13395_ (.CLK(clknet_leaf_124_clk),
    .D(_00614_),
    .Q(\_167_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13396_ (.CLK(clknet_leaf_124_clk),
    .D(_00615_),
    .Q(\_167_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13397_ (.CLK(clknet_leaf_124_clk),
    .D(_00616_),
    .Q(\_167_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13398_ (.CLK(clknet_leaf_125_clk),
    .D(_00617_),
    .Q(\_167_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13399_ (.CLK(clknet_leaf_124_clk),
    .D(_00618_),
    .Q(\_167_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13400_ (.CLK(clknet_leaf_124_clk),
    .D(_00619_),
    .Q(\_167_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13401_ (.CLK(clknet_leaf_125_clk),
    .D(_00620_),
    .Q(\_167_[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13402_ (.CLK(clknet_leaf_130_clk),
    .D(_00621_),
    .Q(\_167_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13403_ (.CLK(clknet_leaf_125_clk),
    .D(_00622_),
    .Q(\_167_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13404_ (.CLK(clknet_leaf_126_clk),
    .D(_00623_),
    .Q(\_167_[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13405_ (.CLK(clknet_leaf_128_clk),
    .D(_00624_),
    .Q(\_167_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13406_ (.CLK(clknet_leaf_126_clk),
    .D(_00625_),
    .Q(\_167_[24] ));
 sky130_fd_sc_hd__dfxtp_2 _13407_ (.CLK(clknet_leaf_127_clk),
    .D(_00626_),
    .Q(\_167_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13408_ (.CLK(clknet_leaf_126_clk),
    .D(_00627_),
    .Q(\_167_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13409_ (.CLK(clknet_leaf_126_clk),
    .D(_00628_),
    .Q(\_167_[27] ));
 sky130_fd_sc_hd__dfxtp_2 _13410_ (.CLK(clknet_leaf_126_clk),
    .D(_00629_),
    .Q(\_167_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13411_ (.CLK(clknet_leaf_126_clk),
    .D(_00630_),
    .Q(\_167_[29] ));
 sky130_fd_sc_hd__dfxtp_2 _13412_ (.CLK(clknet_leaf_128_clk),
    .D(_00631_),
    .Q(\_167_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13413_ (.CLK(clknet_leaf_125_clk),
    .D(_00632_),
    .Q(\_167_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13414_ (.CLK(clknet_leaf_124_clk),
    .D(_00633_),
    .Q(\_164_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13415_ (.CLK(clknet_leaf_12_clk),
    .D(_00634_),
    .Q(\_164_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13416_ (.CLK(clknet_leaf_1_clk),
    .D(_00635_),
    .Q(\_164_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13417_ (.CLK(clknet_leaf_1_clk),
    .D(_00636_),
    .Q(\_164_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13418_ (.CLK(clknet_leaf_3_clk),
    .D(_00637_),
    .Q(\_164_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13419_ (.CLK(clknet_leaf_12_clk),
    .D(_00638_),
    .Q(\_164_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13420_ (.CLK(clknet_leaf_113_clk),
    .D(_00639_),
    .Q(\_164_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13421_ (.CLK(clknet_leaf_1_clk),
    .D(_00640_),
    .Q(\_164_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13422_ (.CLK(clknet_leaf_12_clk),
    .D(_00641_),
    .Q(\_164_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13423_ (.CLK(clknet_leaf_2_clk),
    .D(_00642_),
    .Q(\_164_[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13424_ (.CLK(clknet_leaf_1_clk),
    .D(_00643_),
    .Q(\_164_[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13425_ (.CLK(clknet_leaf_1_clk),
    .D(_00644_),
    .Q(\_164_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13426_ (.CLK(clknet_leaf_113_clk),
    .D(_00645_),
    .Q(\_164_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13427_ (.CLK(clknet_leaf_123_clk),
    .D(_00646_),
    .Q(\_164_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13428_ (.CLK(clknet_leaf_123_clk),
    .D(_00647_),
    .Q(\_164_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13429_ (.CLK(clknet_leaf_123_clk),
    .D(_00648_),
    .Q(\_164_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13430_ (.CLK(clknet_leaf_123_clk),
    .D(_00649_),
    .Q(\_164_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13431_ (.CLK(clknet_leaf_1_clk),
    .D(_00650_),
    .Q(\_164_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13432_ (.CLK(clknet_leaf_123_clk),
    .D(_00651_),
    .Q(\_164_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13433_ (.CLK(clknet_leaf_123_clk),
    .D(_00652_),
    .Q(\_164_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13434_ (.CLK(clknet_leaf_130_clk),
    .D(_00653_),
    .Q(\_164_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13435_ (.CLK(clknet_leaf_125_clk),
    .D(_00654_),
    .Q(\_164_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13436_ (.CLK(clknet_leaf_122_clk),
    .D(_00655_),
    .Q(\_164_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13437_ (.CLK(clknet_leaf_129_clk),
    .D(_00656_),
    .Q(\_164_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13438_ (.CLK(clknet_leaf_126_clk),
    .D(_00657_),
    .Q(\_164_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13439_ (.CLK(clknet_leaf_126_clk),
    .D(_00658_),
    .Q(\_164_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13440_ (.CLK(clknet_leaf_127_clk),
    .D(_00659_),
    .Q(\_164_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13441_ (.CLK(clknet_leaf_122_clk),
    .D(_00660_),
    .Q(\_164_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13442_ (.CLK(clknet_leaf_126_clk),
    .D(_00661_),
    .Q(\_164_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13443_ (.CLK(clknet_leaf_122_clk),
    .D(_00662_),
    .Q(\_164_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13444_ (.CLK(clknet_leaf_128_clk),
    .D(_00663_),
    .Q(\_164_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13445_ (.CLK(clknet_leaf_127_clk),
    .D(_00664_),
    .Q(\_164_[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13446_ (.CLK(clknet_leaf_123_clk),
    .D(_00665_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_4 _13447_ (.CLK(clknet_leaf_12_clk),
    .D(_00666_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_2 _13448_ (.CLK(clknet_leaf_2_clk),
    .D(_00667_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_2 _13449_ (.CLK(clknet_leaf_1_clk),
    .D(_00668_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_2 _13450_ (.CLK(clknet_leaf_3_clk),
    .D(_00669_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_4 _13451_ (.CLK(clknet_leaf_12_clk),
    .D(_00670_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_2 _13452_ (.CLK(clknet_leaf_113_clk),
    .D(_00671_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_4 _13453_ (.CLK(clknet_leaf_2_clk),
    .D(_00672_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_4 _13454_ (.CLK(clknet_leaf_113_clk),
    .D(_00673_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_4 _13455_ (.CLK(clknet_leaf_113_clk),
    .D(_00674_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_4 _13456_ (.CLK(clknet_leaf_1_clk),
    .D(_00675_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_2 _13457_ (.CLK(clknet_leaf_130_clk),
    .D(_00676_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_2 _13458_ (.CLK(clknet_leaf_114_clk),
    .D(_00677_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_2 _13459_ (.CLK(clknet_leaf_123_clk),
    .D(_00678_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_2 _13460_ (.CLK(clknet_leaf_114_clk),
    .D(_00679_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_4 _13461_ (.CLK(clknet_leaf_123_clk),
    .D(_00680_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_4 _13462_ (.CLK(clknet_leaf_123_clk),
    .D(_00681_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_4 _13463_ (.CLK(clknet_leaf_1_clk),
    .D(_00682_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_2 _13464_ (.CLK(clknet_leaf_123_clk),
    .D(_00683_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_2 _13465_ (.CLK(clknet_leaf_123_clk),
    .D(_00684_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_2 _13466_ (.CLK(clknet_leaf_123_clk),
    .D(_00685_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_2 _13467_ (.CLK(clknet_leaf_128_clk),
    .D(_00686_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_4 _13468_ (.CLK(clknet_leaf_122_clk),
    .D(_00687_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _13469_ (.CLK(clknet_leaf_129_clk),
    .D(_00688_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_2 _13470_ (.CLK(clknet_leaf_122_clk),
    .D(_00689_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_4 _13471_ (.CLK(clknet_leaf_122_clk),
    .D(_00690_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_4 _13472_ (.CLK(clknet_leaf_122_clk),
    .D(_00691_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _13473_ (.CLK(clknet_leaf_122_clk),
    .D(_00692_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_4 _13474_ (.CLK(clknet_leaf_127_clk),
    .D(_00693_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_2 _13475_ (.CLK(clknet_leaf_122_clk),
    .D(_00694_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _13476_ (.CLK(clknet_leaf_126_clk),
    .D(_00695_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _13477_ (.CLK(clknet_leaf_127_clk),
    .D(_00696_),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _13478_ (.CLK(clknet_leaf_27_clk),
    .D(_00697_),
    .RESET_B(_00111_),
    .Q(\_190_[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13479_ (.CLK(clknet_leaf_28_clk),
    .D(_00698_),
    .RESET_B(_00112_),
    .Q(\_190_[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13480_ (.CLK(clknet_leaf_28_clk),
    .D(_00699_),
    .RESET_B(_00113_),
    .Q(\_190_[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13481_ (.CLK(clknet_leaf_32_clk),
    .D(_00700_),
    .RESET_B(_00114_),
    .Q(\_190_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13482_ (.CLK(clknet_leaf_35_clk),
    .D(_00701_),
    .Q(\_158_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13483_ (.CLK(clknet_leaf_35_clk),
    .D(_00702_),
    .Q(\_158_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13484_ (.CLK(clknet_leaf_36_clk),
    .D(_00703_),
    .Q(\_158_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13485_ (.CLK(clknet_leaf_36_clk),
    .D(_00704_),
    .Q(\_158_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13486_ (.CLK(clknet_leaf_36_clk),
    .D(_00705_),
    .Q(\_158_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13487_ (.CLK(clknet_leaf_36_clk),
    .D(_00706_),
    .Q(\_158_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13488_ (.CLK(clknet_leaf_50_clk),
    .D(_00707_),
    .Q(\_158_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13489_ (.CLK(clknet_leaf_42_clk),
    .D(_00708_),
    .Q(\_158_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13490_ (.CLK(clknet_leaf_42_clk),
    .D(_00709_),
    .Q(\_158_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13491_ (.CLK(clknet_leaf_46_clk),
    .D(_00710_),
    .Q(\_158_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13492_ (.CLK(clknet_leaf_46_clk),
    .D(_00711_),
    .Q(\_158_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13493_ (.CLK(clknet_leaf_46_clk),
    .D(_00712_),
    .Q(\_158_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13494_ (.CLK(clknet_leaf_41_clk),
    .D(_00713_),
    .Q(\_158_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13495_ (.CLK(clknet_leaf_41_clk),
    .D(_00714_),
    .Q(\_158_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13496_ (.CLK(clknet_leaf_41_clk),
    .D(_00715_),
    .Q(\_158_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13497_ (.CLK(clknet_leaf_41_clk),
    .D(_00716_),
    .Q(\_158_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13498_ (.CLK(clknet_leaf_50_clk),
    .D(_00717_),
    .Q(\_158_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13499_ (.CLK(clknet_leaf_36_clk),
    .D(_00718_),
    .Q(\_158_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13500_ (.CLK(clknet_leaf_36_clk),
    .D(_00719_),
    .Q(\_158_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13501_ (.CLK(clknet_leaf_36_clk),
    .D(_00720_),
    .Q(\_158_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13502_ (.CLK(clknet_leaf_37_clk),
    .D(_00721_),
    .Q(\_158_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13503_ (.CLK(clknet_leaf_37_clk),
    .D(_00722_),
    .Q(\_158_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13504_ (.CLK(clknet_leaf_56_clk),
    .D(_00723_),
    .Q(\_152_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13505_ (.CLK(clknet_leaf_57_clk),
    .D(_00724_),
    .Q(\_152_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13506_ (.CLK(clknet_leaf_60_clk),
    .D(_00725_),
    .Q(\_152_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13507_ (.CLK(clknet_leaf_60_clk),
    .D(_00726_),
    .Q(\_152_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13508_ (.CLK(clknet_leaf_58_clk),
    .D(_00727_),
    .Q(\_152_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13509_ (.CLK(clknet_leaf_60_clk),
    .D(_00728_),
    .Q(\_152_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13510_ (.CLK(clknet_leaf_60_clk),
    .D(_00729_),
    .Q(\_152_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13511_ (.CLK(clknet_leaf_60_clk),
    .D(_00730_),
    .Q(\_152_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13512_ (.CLK(clknet_leaf_55_clk),
    .D(_00731_),
    .Q(\_152_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13513_ (.CLK(clknet_leaf_55_clk),
    .D(_00732_),
    .Q(\_152_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13514_ (.CLK(clknet_leaf_55_clk),
    .D(_00733_),
    .Q(\_152_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13515_ (.CLK(clknet_leaf_81_clk),
    .D(_00734_),
    .Q(\_152_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13516_ (.CLK(clknet_leaf_78_clk),
    .D(_00735_),
    .Q(\_152_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13517_ (.CLK(clknet_leaf_80_clk),
    .D(_00736_),
    .Q(\_152_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13518_ (.CLK(clknet_leaf_81_clk),
    .D(_00737_),
    .Q(\_152_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13519_ (.CLK(clknet_leaf_78_clk),
    .D(_00738_),
    .Q(\_152_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13520_ (.CLK(clknet_leaf_79_clk),
    .D(_00739_),
    .Q(\_152_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13521_ (.CLK(clknet_leaf_81_clk),
    .D(_00740_),
    .Q(\_152_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13522_ (.CLK(clknet_leaf_80_clk),
    .D(_00741_),
    .Q(\_152_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13523_ (.CLK(clknet_leaf_78_clk),
    .D(_00742_),
    .Q(\_152_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13524_ (.CLK(clknet_leaf_75_clk),
    .D(_00743_),
    .Q(\_152_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13525_ (.CLK(clknet_leaf_78_clk),
    .D(_00744_),
    .Q(\_152_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13526_ (.CLK(clknet_leaf_76_clk),
    .D(_00745_),
    .Q(\_152_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13527_ (.CLK(clknet_leaf_76_clk),
    .D(_00746_),
    .Q(\_152_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13528_ (.CLK(clknet_leaf_47_clk),
    .D(_00747_),
    .Q(\_152_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13529_ (.CLK(clknet_leaf_47_clk),
    .D(_00748_),
    .Q(\_152_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13530_ (.CLK(clknet_leaf_67_clk),
    .D(_00749_),
    .Q(\_152_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13531_ (.CLK(clknet_leaf_67_clk),
    .D(_00750_),
    .Q(\_152_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13532_ (.CLK(clknet_leaf_67_clk),
    .D(_00751_),
    .Q(\_152_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13533_ (.CLK(clknet_leaf_67_clk),
    .D(_00752_),
    .Q(\_152_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13534_ (.CLK(clknet_leaf_66_clk),
    .D(_00753_),
    .Q(\_152_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13535_ (.CLK(clknet_leaf_66_clk),
    .D(_00754_),
    .Q(\_152_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13536_ (.CLK(clknet_leaf_68_clk),
    .D(_00755_),
    .Q(\_149_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13537_ (.CLK(clknet_leaf_66_clk),
    .D(_00756_),
    .Q(\_149_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13538_ (.CLK(clknet_leaf_66_clk),
    .D(_00757_),
    .Q(\_149_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13539_ (.CLK(clknet_leaf_65_clk),
    .D(_00758_),
    .Q(\_149_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13540_ (.CLK(clknet_leaf_65_clk),
    .D(_00759_),
    .Q(\_149_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13541_ (.CLK(clknet_leaf_63_clk),
    .D(_00760_),
    .Q(\_149_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13542_ (.CLK(clknet_leaf_65_clk),
    .D(_00761_),
    .Q(\_149_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13543_ (.CLK(clknet_leaf_73_clk),
    .D(_00762_),
    .Q(\_149_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13544_ (.CLK(clknet_leaf_74_clk),
    .D(_00763_),
    .Q(\_149_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13545_ (.CLK(clknet_leaf_68_clk),
    .D(_00764_),
    .Q(\_149_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13546_ (.CLK(clknet_leaf_87_clk),
    .D(_00765_),
    .Q(\_149_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13547_ (.CLK(clknet_leaf_84_clk),
    .D(_00766_),
    .Q(\_149_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13548_ (.CLK(clknet_leaf_84_clk),
    .D(_00767_),
    .Q(\_149_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13549_ (.CLK(clknet_leaf_87_clk),
    .D(_00768_),
    .Q(\_149_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13550_ (.CLK(clknet_leaf_86_clk),
    .D(_00769_),
    .Q(\_149_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13551_ (.CLK(clknet_leaf_87_clk),
    .D(_00770_),
    .Q(\_149_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13552_ (.CLK(clknet_leaf_84_clk),
    .D(_00771_),
    .Q(\_149_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13553_ (.CLK(clknet_leaf_79_clk),
    .D(_00772_),
    .Q(\_149_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13554_ (.CLK(clknet_leaf_74_clk),
    .D(_00773_),
    .Q(\_149_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13555_ (.CLK(clknet_leaf_74_clk),
    .D(_00774_),
    .Q(\_149_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13556_ (.CLK(clknet_leaf_73_clk),
    .D(_00775_),
    .Q(\_149_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13557_ (.CLK(clknet_leaf_73_clk),
    .D(_00776_),
    .Q(\_149_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13558_ (.CLK(clknet_leaf_76_clk),
    .D(_00777_),
    .Q(\_149_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13559_ (.CLK(clknet_leaf_75_clk),
    .D(_00778_),
    .Q(\_149_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13560_ (.CLK(clknet_leaf_74_clk),
    .D(_00779_),
    .Q(\_149_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13561_ (.CLK(clknet_leaf_75_clk),
    .D(_00780_),
    .Q(\_149_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13562_ (.CLK(clknet_leaf_75_clk),
    .D(_00781_),
    .Q(\_149_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13563_ (.CLK(clknet_leaf_75_clk),
    .D(_00782_),
    .Q(\_149_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13564_ (.CLK(clknet_leaf_75_clk),
    .D(_00783_),
    .Q(\_149_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13565_ (.CLK(clknet_leaf_76_clk),
    .D(_00784_),
    .Q(\_149_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13566_ (.CLK(clknet_leaf_75_clk),
    .D(_00785_),
    .Q(\_149_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13567_ (.CLK(clknet_leaf_68_clk),
    .D(_00786_),
    .Q(\_149_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13568_ (.CLK(clknet_leaf_55_clk),
    .D(_00787_),
    .Q(\_142_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13569_ (.CLK(clknet_leaf_54_clk),
    .D(_00788_),
    .Q(\_142_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13570_ (.CLK(clknet_leaf_34_clk),
    .D(_00789_),
    .Q(\_142_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13571_ (.CLK(clknet_leaf_34_clk),
    .D(_00790_),
    .Q(\_142_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13572_ (.CLK(clknet_leaf_52_clk),
    .D(_00791_),
    .Q(\_142_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13573_ (.CLK(clknet_leaf_53_clk),
    .D(_00792_),
    .Q(\_142_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13574_ (.CLK(clknet_leaf_34_clk),
    .D(_00793_),
    .Q(\_142_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13575_ (.CLK(clknet_leaf_54_clk),
    .D(_00794_),
    .Q(\_142_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13576_ (.CLK(clknet_leaf_54_clk),
    .D(_00795_),
    .Q(\_142_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13577_ (.CLK(clknet_leaf_52_clk),
    .D(_00796_),
    .Q(\_142_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13578_ (.CLK(clknet_leaf_35_clk),
    .D(_00797_),
    .Q(\_142_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13579_ (.CLK(clknet_leaf_51_clk),
    .D(_00798_),
    .Q(\_142_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13580_ (.CLK(clknet_leaf_51_clk),
    .D(_00799_),
    .Q(\_142_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13581_ (.CLK(clknet_leaf_51_clk),
    .D(_00800_),
    .Q(\_142_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13582_ (.CLK(clknet_leaf_45_clk),
    .D(_00801_),
    .Q(\_142_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13583_ (.CLK(clknet_leaf_45_clk),
    .D(_00802_),
    .Q(\_142_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13584_ (.CLK(clknet_leaf_45_clk),
    .D(_00803_),
    .Q(\_142_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13585_ (.CLK(clknet_leaf_45_clk),
    .D(_00804_),
    .Q(\_142_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13586_ (.CLK(clknet_leaf_46_clk),
    .D(_00805_),
    .Q(\_142_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13587_ (.CLK(clknet_leaf_46_clk),
    .D(_00806_),
    .Q(\_142_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13588_ (.CLK(clknet_leaf_46_clk),
    .D(_00807_),
    .Q(\_142_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13589_ (.CLK(clknet_leaf_50_clk),
    .D(_00808_),
    .Q(\_142_[21] ));
 sky130_fd_sc_hd__dfxtp_2 _13590_ (.CLK(clknet_leaf_48_clk),
    .D(_00809_),
    .Q(\_142_[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13591_ (.CLK(clknet_leaf_46_clk),
    .D(_00810_),
    .Q(\_142_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13592_ (.CLK(clknet_leaf_50_clk),
    .D(_00811_),
    .Q(\_142_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13593_ (.CLK(clknet_leaf_49_clk),
    .D(_00812_),
    .Q(\_142_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13594_ (.CLK(clknet_leaf_49_clk),
    .D(_00813_),
    .Q(\_142_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13595_ (.CLK(clknet_leaf_50_clk),
    .D(_00814_),
    .Q(\_142_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13596_ (.CLK(clknet_leaf_50_clk),
    .D(_00815_),
    .Q(\_142_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13597_ (.CLK(clknet_leaf_36_clk),
    .D(_00816_),
    .Q(\_142_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13598_ (.CLK(clknet_leaf_51_clk),
    .D(_00817_),
    .Q(\_142_[30] ));
 sky130_fd_sc_hd__dfxtp_2 _13599_ (.CLK(clknet_leaf_56_clk),
    .D(_00818_),
    .Q(\_142_[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13600_ (.CLK(clknet_leaf_53_clk),
    .D(_00819_),
    .Q(\_140_[0] ));
 sky130_fd_sc_hd__dfxtp_2 _13601_ (.CLK(clknet_leaf_53_clk),
    .D(_00820_),
    .Q(\_140_[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13602_ (.CLK(clknet_leaf_52_clk),
    .D(_00821_),
    .Q(\_140_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13603_ (.CLK(clknet_leaf_52_clk),
    .D(_00822_),
    .Q(\_140_[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13604_ (.CLK(clknet_leaf_52_clk),
    .D(_00823_),
    .Q(\_140_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13605_ (.CLK(clknet_leaf_53_clk),
    .D(_00824_),
    .Q(\_140_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13606_ (.CLK(clknet_leaf_52_clk),
    .D(_00825_),
    .Q(\_140_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13607_ (.CLK(clknet_leaf_53_clk),
    .D(_00826_),
    .Q(\_140_[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13608_ (.CLK(clknet_leaf_53_clk),
    .D(_00827_),
    .Q(\_140_[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13609_ (.CLK(clknet_leaf_52_clk),
    .D(_00828_),
    .Q(\_140_[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13610_ (.CLK(clknet_leaf_52_clk),
    .D(_00829_),
    .Q(\_140_[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13611_ (.CLK(clknet_leaf_52_clk),
    .D(_00830_),
    .Q(\_140_[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13612_ (.CLK(clknet_leaf_51_clk),
    .D(_00831_),
    .Q(\_140_[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13613_ (.CLK(clknet_leaf_51_clk),
    .D(_00832_),
    .Q(\_140_[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13614_ (.CLK(clknet_leaf_49_clk),
    .D(_00833_),
    .Q(\_140_[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13615_ (.CLK(clknet_leaf_45_clk),
    .D(_00834_),
    .Q(\_140_[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13616_ (.CLK(clknet_leaf_47_clk),
    .D(_00835_),
    .Q(\_140_[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13617_ (.CLK(clknet_leaf_45_clk),
    .D(_00836_),
    .Q(\_140_[17] ));
 sky130_fd_sc_hd__dfxtp_2 _13618_ (.CLK(clknet_leaf_49_clk),
    .D(_00837_),
    .Q(\_140_[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13619_ (.CLK(clknet_leaf_46_clk),
    .D(_00838_),
    .Q(\_140_[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13620_ (.CLK(clknet_leaf_46_clk),
    .D(_00839_),
    .Q(\_140_[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13621_ (.CLK(clknet_leaf_49_clk),
    .D(_00840_),
    .Q(\_140_[21] ));
 sky130_fd_sc_hd__dfxtp_2 _13622_ (.CLK(clknet_leaf_49_clk),
    .D(_00841_),
    .Q(\_140_[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13623_ (.CLK(clknet_leaf_50_clk),
    .D(_00842_),
    .Q(\_140_[23] ));
 sky130_fd_sc_hd__dfxtp_2 _13624_ (.CLK(clknet_leaf_50_clk),
    .D(_00843_),
    .Q(\_140_[24] ));
 sky130_fd_sc_hd__dfxtp_2 _13625_ (.CLK(clknet_leaf_49_clk),
    .D(_00844_),
    .Q(\_140_[25] ));
 sky130_fd_sc_hd__dfxtp_2 _13626_ (.CLK(clknet_leaf_51_clk),
    .D(_00845_),
    .Q(\_140_[26] ));
 sky130_fd_sc_hd__dfxtp_2 _13627_ (.CLK(clknet_leaf_50_clk),
    .D(_00846_),
    .Q(\_140_[27] ));
 sky130_fd_sc_hd__dfxtp_2 _13628_ (.CLK(clknet_leaf_51_clk),
    .D(_00847_),
    .Q(\_140_[28] ));
 sky130_fd_sc_hd__dfxtp_2 _13629_ (.CLK(clknet_leaf_51_clk),
    .D(_00848_),
    .Q(\_140_[29] ));
 sky130_fd_sc_hd__dfxtp_2 _13630_ (.CLK(clknet_leaf_51_clk),
    .D(_00849_),
    .Q(\_140_[30] ));
 sky130_fd_sc_hd__dfxtp_2 _13631_ (.CLK(clknet_leaf_53_clk),
    .D(_00850_),
    .Q(\_140_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13632_ (.CLK(clknet_leaf_58_clk),
    .D(_00851_),
    .Q(\_138_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13633_ (.CLK(clknet_leaf_58_clk),
    .D(_00852_),
    .Q(\_138_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13634_ (.CLK(clknet_leaf_54_clk),
    .D(_00853_),
    .Q(\_138_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13635_ (.CLK(clknet_leaf_53_clk),
    .D(_00854_),
    .Q(\_138_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13636_ (.CLK(clknet_leaf_53_clk),
    .D(_00855_),
    .Q(\_138_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13637_ (.CLK(clknet_leaf_54_clk),
    .D(_00856_),
    .Q(\_138_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13638_ (.CLK(clknet_leaf_53_clk),
    .D(_00857_),
    .Q(\_138_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13639_ (.CLK(clknet_leaf_53_clk),
    .D(_00858_),
    .Q(\_138_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13640_ (.CLK(clknet_leaf_54_clk),
    .D(_00859_),
    .Q(\_138_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13641_ (.CLK(clknet_leaf_54_clk),
    .D(_00860_),
    .Q(\_138_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13642_ (.CLK(clknet_leaf_48_clk),
    .D(_00861_),
    .Q(\_138_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13643_ (.CLK(clknet_leaf_48_clk),
    .D(_00862_),
    .Q(\_138_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13644_ (.CLK(clknet_leaf_78_clk),
    .D(_00863_),
    .Q(\_138_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13645_ (.CLK(clknet_leaf_47_clk),
    .D(_00864_),
    .Q(\_138_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13646_ (.CLK(clknet_leaf_47_clk),
    .D(_00865_),
    .Q(\_138_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13647_ (.CLK(clknet_leaf_47_clk),
    .D(_00866_),
    .Q(\_138_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13648_ (.CLK(clknet_leaf_47_clk),
    .D(_00867_),
    .Q(\_138_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13649_ (.CLK(clknet_leaf_78_clk),
    .D(_00868_),
    .Q(\_138_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13650_ (.CLK(clknet_leaf_47_clk),
    .D(_00869_),
    .Q(\_138_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13651_ (.CLK(clknet_leaf_77_clk),
    .D(_00870_),
    .Q(\_138_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13652_ (.CLK(clknet_leaf_48_clk),
    .D(_00871_),
    .Q(\_138_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13653_ (.CLK(clknet_leaf_47_clk),
    .D(_00872_),
    .Q(\_138_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13654_ (.CLK(clknet_leaf_56_clk),
    .D(_00873_),
    .Q(\_138_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13655_ (.CLK(clknet_leaf_48_clk),
    .D(_00874_),
    .Q(\_138_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13656_ (.CLK(clknet_leaf_56_clk),
    .D(_00875_),
    .Q(\_138_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13657_ (.CLK(clknet_leaf_56_clk),
    .D(_00876_),
    .Q(\_138_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13658_ (.CLK(clknet_leaf_56_clk),
    .D(_00877_),
    .Q(\_138_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13659_ (.CLK(clknet_leaf_56_clk),
    .D(_00878_),
    .Q(\_138_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13660_ (.CLK(clknet_leaf_56_clk),
    .D(_00879_),
    .Q(\_138_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13661_ (.CLK(clknet_leaf_56_clk),
    .D(_00880_),
    .Q(\_138_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13662_ (.CLK(clknet_leaf_58_clk),
    .D(_00881_),
    .Q(\_138_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13663_ (.CLK(clknet_leaf_55_clk),
    .D(_00882_),
    .Q(\_138_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13664_ (.CLK(clknet_leaf_58_clk),
    .D(_00883_),
    .Q(\_136_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13665_ (.CLK(clknet_leaf_59_clk),
    .D(_00884_),
    .Q(\_136_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13666_ (.CLK(clknet_leaf_54_clk),
    .D(_00885_),
    .Q(\_136_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13667_ (.CLK(clknet_leaf_59_clk),
    .D(_00886_),
    .Q(\_136_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13668_ (.CLK(clknet_leaf_54_clk),
    .D(_00887_),
    .Q(\_136_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13669_ (.CLK(clknet_leaf_59_clk),
    .D(_00888_),
    .Q(\_136_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13670_ (.CLK(clknet_leaf_54_clk),
    .D(_00889_),
    .Q(\_136_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13671_ (.CLK(clknet_leaf_54_clk),
    .D(_00890_),
    .Q(\_136_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13672_ (.CLK(clknet_leaf_54_clk),
    .D(_00891_),
    .Q(\_136_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13673_ (.CLK(clknet_leaf_54_clk),
    .D(_00892_),
    .Q(\_136_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13674_ (.CLK(clknet_leaf_48_clk),
    .D(_00893_),
    .Q(\_136_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13675_ (.CLK(clknet_leaf_48_clk),
    .D(_00894_),
    .Q(\_136_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13676_ (.CLK(clknet_leaf_77_clk),
    .D(_00895_),
    .Q(\_136_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13677_ (.CLK(clknet_leaf_78_clk),
    .D(_00896_),
    .Q(\_136_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13678_ (.CLK(clknet_leaf_47_clk),
    .D(_00897_),
    .Q(\_136_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13679_ (.CLK(clknet_leaf_78_clk),
    .D(_00898_),
    .Q(\_136_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13680_ (.CLK(clknet_leaf_78_clk),
    .D(_00899_),
    .Q(\_136_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13681_ (.CLK(clknet_leaf_78_clk),
    .D(_00900_),
    .Q(\_136_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13682_ (.CLK(clknet_leaf_77_clk),
    .D(_00901_),
    .Q(\_136_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13683_ (.CLK(clknet_leaf_77_clk),
    .D(_00902_),
    .Q(\_136_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13684_ (.CLK(clknet_leaf_77_clk),
    .D(_00903_),
    .Q(\_136_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13685_ (.CLK(clknet_leaf_77_clk),
    .D(_00904_),
    .Q(\_136_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13686_ (.CLK(clknet_leaf_56_clk),
    .D(_00905_),
    .Q(\_136_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13687_ (.CLK(clknet_leaf_67_clk),
    .D(_00906_),
    .Q(\_136_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13688_ (.CLK(clknet_leaf_56_clk),
    .D(_00907_),
    .Q(\_136_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13689_ (.CLK(clknet_leaf_56_clk),
    .D(_00908_),
    .Q(\_136_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13690_ (.CLK(clknet_leaf_56_clk),
    .D(_00909_),
    .Q(\_136_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13691_ (.CLK(clknet_leaf_57_clk),
    .D(_00910_),
    .Q(\_136_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13692_ (.CLK(clknet_leaf_57_clk),
    .D(_00911_),
    .Q(\_136_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13693_ (.CLK(clknet_leaf_57_clk),
    .D(_00912_),
    .Q(\_136_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13694_ (.CLK(clknet_leaf_58_clk),
    .D(_00913_),
    .Q(\_136_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13695_ (.CLK(clknet_leaf_58_clk),
    .D(_00914_),
    .Q(\_136_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13696_ (.CLK(clknet_leaf_59_clk),
    .D(_00915_),
    .Q(\_134_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13697_ (.CLK(clknet_leaf_59_clk),
    .D(_00916_),
    .Q(\_134_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13698_ (.CLK(clknet_leaf_59_clk),
    .D(_00917_),
    .Q(\_134_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13699_ (.CLK(clknet_leaf_59_clk),
    .D(_00918_),
    .Q(\_134_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13700_ (.CLK(clknet_leaf_58_clk),
    .D(_00919_),
    .Q(\_134_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13701_ (.CLK(clknet_leaf_59_clk),
    .D(_00920_),
    .Q(\_134_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13702_ (.CLK(clknet_leaf_59_clk),
    .D(_00921_),
    .Q(\_134_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13703_ (.CLK(clknet_leaf_59_clk),
    .D(_00922_),
    .Q(\_134_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13704_ (.CLK(clknet_leaf_54_clk),
    .D(_00923_),
    .Q(\_134_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13705_ (.CLK(clknet_leaf_55_clk),
    .D(_00924_),
    .Q(\_134_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13706_ (.CLK(clknet_leaf_48_clk),
    .D(_00925_),
    .Q(\_134_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13707_ (.CLK(clknet_leaf_48_clk),
    .D(_00926_),
    .Q(\_134_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13708_ (.CLK(clknet_leaf_77_clk),
    .D(_00927_),
    .Q(\_134_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13709_ (.CLK(clknet_leaf_78_clk),
    .D(_00928_),
    .Q(\_134_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13710_ (.CLK(clknet_leaf_78_clk),
    .D(_00929_),
    .Q(\_134_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13711_ (.CLK(clknet_leaf_78_clk),
    .D(_00930_),
    .Q(\_134_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13712_ (.CLK(clknet_leaf_78_clk),
    .D(_00931_),
    .Q(\_134_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13713_ (.CLK(clknet_leaf_77_clk),
    .D(_00932_),
    .Q(\_134_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13714_ (.CLK(clknet_leaf_77_clk),
    .D(_00933_),
    .Q(\_134_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13715_ (.CLK(clknet_leaf_77_clk),
    .D(_00934_),
    .Q(\_134_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13716_ (.CLK(clknet_leaf_77_clk),
    .D(_00935_),
    .Q(\_134_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13717_ (.CLK(clknet_leaf_77_clk),
    .D(_00936_),
    .Q(\_134_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13718_ (.CLK(clknet_leaf_67_clk),
    .D(_00937_),
    .Q(\_134_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13719_ (.CLK(clknet_leaf_67_clk),
    .D(_00938_),
    .Q(\_134_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13720_ (.CLK(clknet_leaf_67_clk),
    .D(_00939_),
    .Q(\_134_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13721_ (.CLK(clknet_leaf_56_clk),
    .D(_00940_),
    .Q(\_134_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13722_ (.CLK(clknet_leaf_57_clk),
    .D(_00941_),
    .Q(\_134_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13723_ (.CLK(clknet_leaf_57_clk),
    .D(_00942_),
    .Q(\_134_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13724_ (.CLK(clknet_leaf_57_clk),
    .D(_00943_),
    .Q(\_134_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13725_ (.CLK(clknet_leaf_57_clk),
    .D(_00944_),
    .Q(\_134_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13726_ (.CLK(clknet_leaf_57_clk),
    .D(_00945_),
    .Q(\_134_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13727_ (.CLK(clknet_leaf_58_clk),
    .D(_00946_),
    .Q(\_134_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13728_ (.CLK(clknet_leaf_66_clk),
    .D(_00947_),
    .Q(\_132_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13729_ (.CLK(clknet_leaf_57_clk),
    .D(_00948_),
    .Q(\_132_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13730_ (.CLK(clknet_leaf_59_clk),
    .D(_00949_),
    .Q(\_132_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13731_ (.CLK(clknet_leaf_60_clk),
    .D(_00950_),
    .Q(\_132_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13732_ (.CLK(clknet_leaf_60_clk),
    .D(_00951_),
    .Q(\_132_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13733_ (.CLK(clknet_leaf_61_clk),
    .D(_00952_),
    .Q(\_132_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13734_ (.CLK(clknet_leaf_59_clk),
    .D(_00953_),
    .Q(\_132_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13735_ (.CLK(clknet_leaf_59_clk),
    .D(_00954_),
    .Q(\_132_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13736_ (.CLK(clknet_leaf_55_clk),
    .D(_00955_),
    .Q(\_132_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13737_ (.CLK(clknet_leaf_58_clk),
    .D(_00956_),
    .Q(\_132_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13738_ (.CLK(clknet_leaf_77_clk),
    .D(_00957_),
    .Q(\_132_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13739_ (.CLK(clknet_leaf_48_clk),
    .D(_00958_),
    .Q(\_132_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13740_ (.CLK(clknet_leaf_78_clk),
    .D(_00959_),
    .Q(\_132_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13741_ (.CLK(clknet_leaf_80_clk),
    .D(_00960_),
    .Q(\_132_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13742_ (.CLK(clknet_leaf_78_clk),
    .D(_00961_),
    .Q(\_132_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13743_ (.CLK(clknet_leaf_79_clk),
    .D(_00962_),
    .Q(\_132_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13744_ (.CLK(clknet_leaf_79_clk),
    .D(_00963_),
    .Q(\_132_[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13745_ (.CLK(clknet_leaf_79_clk),
    .D(_00964_),
    .Q(\_132_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13746_ (.CLK(clknet_leaf_74_clk),
    .D(_00965_),
    .Q(\_132_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13747_ (.CLK(clknet_leaf_74_clk),
    .D(_00966_),
    .Q(\_132_[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13748_ (.CLK(clknet_leaf_77_clk),
    .D(_00967_),
    .Q(\_132_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13749_ (.CLK(clknet_leaf_75_clk),
    .D(_00968_),
    .Q(\_132_[21] ));
 sky130_fd_sc_hd__dfxtp_2 _13750_ (.CLK(clknet_leaf_67_clk),
    .D(_00969_),
    .Q(\_132_[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13751_ (.CLK(clknet_leaf_67_clk),
    .D(_00970_),
    .Q(\_132_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13752_ (.CLK(clknet_leaf_67_clk),
    .D(_00971_),
    .Q(\_132_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13753_ (.CLK(clknet_leaf_67_clk),
    .D(_00972_),
    .Q(\_132_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13754_ (.CLK(clknet_leaf_66_clk),
    .D(_00973_),
    .Q(\_132_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13755_ (.CLK(clknet_leaf_57_clk),
    .D(_00974_),
    .Q(\_132_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13756_ (.CLK(clknet_leaf_67_clk),
    .D(_00975_),
    .Q(\_132_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13757_ (.CLK(clknet_leaf_57_clk),
    .D(_00976_),
    .Q(\_132_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13758_ (.CLK(clknet_leaf_57_clk),
    .D(_00977_),
    .Q(\_132_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13759_ (.CLK(clknet_leaf_57_clk),
    .D(_00978_),
    .Q(\_132_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13760_ (.CLK(clknet_leaf_65_clk),
    .D(_00979_),
    .Q(\_130_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13761_ (.CLK(clknet_leaf_66_clk),
    .D(_00980_),
    .Q(\_130_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13762_ (.CLK(clknet_leaf_63_clk),
    .D(_00981_),
    .Q(\_130_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13763_ (.CLK(clknet_leaf_63_clk),
    .D(_00982_),
    .Q(\_130_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13764_ (.CLK(clknet_leaf_62_clk),
    .D(_00983_),
    .Q(\_130_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13765_ (.CLK(clknet_leaf_62_clk),
    .D(_00984_),
    .Q(\_130_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13766_ (.CLK(clknet_leaf_60_clk),
    .D(_00985_),
    .Q(\_130_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13767_ (.CLK(clknet_leaf_60_clk),
    .D(_00986_),
    .Q(\_130_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13768_ (.CLK(clknet_leaf_58_clk),
    .D(_00987_),
    .Q(\_130_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13769_ (.CLK(clknet_leaf_58_clk),
    .D(_00988_),
    .Q(\_130_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13770_ (.CLK(clknet_leaf_87_clk),
    .D(_00989_),
    .Q(\_130_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13771_ (.CLK(clknet_leaf_87_clk),
    .D(_00990_),
    .Q(\_130_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13772_ (.CLK(clknet_leaf_87_clk),
    .D(_00991_),
    .Q(\_130_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13773_ (.CLK(clknet_leaf_84_clk),
    .D(_00992_),
    .Q(\_130_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13774_ (.CLK(clknet_leaf_84_clk),
    .D(_00993_),
    .Q(\_130_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13775_ (.CLK(clknet_leaf_84_clk),
    .D(_00994_),
    .Q(\_130_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13776_ (.CLK(clknet_leaf_93_clk),
    .D(_00995_),
    .Q(\_130_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13777_ (.CLK(clknet_leaf_95_clk),
    .D(_00996_),
    .Q(\_130_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13778_ (.CLK(clknet_leaf_94_clk),
    .D(_00997_),
    .Q(\_130_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13779_ (.CLK(clknet_leaf_94_clk),
    .D(_00998_),
    .Q(\_130_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13780_ (.CLK(clknet_leaf_93_clk),
    .D(_00999_),
    .Q(\_130_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13781_ (.CLK(clknet_leaf_93_clk),
    .D(_01000_),
    .Q(\_130_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13782_ (.CLK(clknet_leaf_94_clk),
    .D(_01001_),
    .Q(\_130_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13783_ (.CLK(clknet_leaf_94_clk),
    .D(_01002_),
    .Q(\_130_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13784_ (.CLK(clknet_leaf_76_clk),
    .D(_01003_),
    .Q(\_130_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13785_ (.CLK(clknet_leaf_76_clk),
    .D(_01004_),
    .Q(\_130_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13786_ (.CLK(clknet_leaf_68_clk),
    .D(_01005_),
    .Q(\_130_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13787_ (.CLK(clknet_leaf_68_clk),
    .D(_01006_),
    .Q(\_130_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13788_ (.CLK(clknet_leaf_68_clk),
    .D(_01007_),
    .Q(\_130_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13789_ (.CLK(clknet_leaf_69_clk),
    .D(_01008_),
    .Q(\_130_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13790_ (.CLK(clknet_leaf_65_clk),
    .D(_01009_),
    .Q(\_130_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13791_ (.CLK(clknet_leaf_65_clk),
    .D(_01010_),
    .Q(\_130_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13792_ (.CLK(clknet_leaf_65_clk),
    .D(_01011_),
    .Q(\_128_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13793_ (.CLK(clknet_leaf_63_clk),
    .D(_01012_),
    .Q(\_128_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13794_ (.CLK(clknet_leaf_63_clk),
    .D(_01013_),
    .Q(\_128_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13795_ (.CLK(clknet_leaf_63_clk),
    .D(_01014_),
    .Q(\_128_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13796_ (.CLK(clknet_leaf_62_clk),
    .D(_01015_),
    .Q(\_128_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13797_ (.CLK(clknet_leaf_63_clk),
    .D(_01016_),
    .Q(\_128_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13798_ (.CLK(clknet_leaf_60_clk),
    .D(_01017_),
    .Q(\_128_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13799_ (.CLK(clknet_leaf_61_clk),
    .D(_01018_),
    .Q(\_128_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13800_ (.CLK(clknet_leaf_58_clk),
    .D(_01019_),
    .Q(\_128_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13801_ (.CLK(clknet_leaf_60_clk),
    .D(_01020_),
    .Q(\_128_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13802_ (.CLK(clknet_leaf_86_clk),
    .D(_01021_),
    .Q(\_128_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13803_ (.CLK(clknet_leaf_93_clk),
    .D(_01022_),
    .Q(\_128_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13804_ (.CLK(clknet_leaf_87_clk),
    .D(_01023_),
    .Q(\_128_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13805_ (.CLK(clknet_leaf_93_clk),
    .D(_01024_),
    .Q(\_128_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13806_ (.CLK(clknet_leaf_98_clk),
    .D(_01025_),
    .Q(\_128_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13807_ (.CLK(clknet_leaf_98_clk),
    .D(_01026_),
    .Q(\_128_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13808_ (.CLK(clknet_leaf_95_clk),
    .D(_01027_),
    .Q(\_128_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13809_ (.CLK(clknet_leaf_95_clk),
    .D(_01028_),
    .Q(\_128_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13810_ (.CLK(clknet_leaf_94_clk),
    .D(_01029_),
    .Q(\_128_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13811_ (.CLK(clknet_leaf_95_clk),
    .D(_01030_),
    .Q(\_128_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13812_ (.CLK(clknet_leaf_94_clk),
    .D(_01031_),
    .Q(\_128_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13813_ (.CLK(clknet_leaf_93_clk),
    .D(_01032_),
    .Q(\_128_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13814_ (.CLK(clknet_leaf_94_clk),
    .D(_01033_),
    .Q(\_128_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13815_ (.CLK(clknet_leaf_93_clk),
    .D(_01034_),
    .Q(\_128_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13816_ (.CLK(clknet_leaf_68_clk),
    .D(_01035_),
    .Q(\_128_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13817_ (.CLK(clknet_leaf_71_clk),
    .D(_01036_),
    .Q(\_128_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13818_ (.CLK(clknet_leaf_75_clk),
    .D(_01037_),
    .Q(\_128_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13819_ (.CLK(clknet_leaf_71_clk),
    .D(_01038_),
    .Q(\_128_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13820_ (.CLK(clknet_leaf_68_clk),
    .D(_01039_),
    .Q(\_128_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13821_ (.CLK(clknet_leaf_68_clk),
    .D(_01040_),
    .Q(\_128_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13822_ (.CLK(clknet_leaf_69_clk),
    .D(_01041_),
    .Q(\_128_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13823_ (.CLK(clknet_leaf_65_clk),
    .D(_01042_),
    .Q(\_128_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13824_ (.CLK(clknet_leaf_64_clk),
    .D(_01043_),
    .Q(\_126_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13825_ (.CLK(clknet_leaf_64_clk),
    .D(_01044_),
    .Q(\_126_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13826_ (.CLK(clknet_leaf_63_clk),
    .D(_01045_),
    .Q(\_126_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13827_ (.CLK(clknet_leaf_63_clk),
    .D(_01046_),
    .Q(\_126_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13828_ (.CLK(clknet_leaf_63_clk),
    .D(_01047_),
    .Q(\_126_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13829_ (.CLK(clknet_leaf_63_clk),
    .D(_01048_),
    .Q(\_126_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13830_ (.CLK(clknet_leaf_61_clk),
    .D(_01049_),
    .Q(\_126_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13831_ (.CLK(clknet_leaf_62_clk),
    .D(_01050_),
    .Q(\_126_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13832_ (.CLK(clknet_leaf_62_clk),
    .D(_01051_),
    .Q(\_126_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13833_ (.CLK(clknet_leaf_62_clk),
    .D(_01052_),
    .Q(\_126_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13834_ (.CLK(clknet_leaf_93_clk),
    .D(_01053_),
    .Q(\_126_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13835_ (.CLK(clknet_leaf_93_clk),
    .D(_01054_),
    .Q(\_126_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13836_ (.CLK(clknet_leaf_98_clk),
    .D(_01055_),
    .Q(\_126_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13837_ (.CLK(clknet_leaf_95_clk),
    .D(_01056_),
    .Q(\_126_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13838_ (.CLK(clknet_leaf_98_clk),
    .D(_01057_),
    .Q(\_126_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13839_ (.CLK(clknet_leaf_95_clk),
    .D(_01058_),
    .Q(\_126_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13840_ (.CLK(clknet_leaf_95_clk),
    .D(_01059_),
    .Q(\_126_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13841_ (.CLK(clknet_leaf_95_clk),
    .D(_01060_),
    .Q(\_126_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13842_ (.CLK(clknet_leaf_94_clk),
    .D(_01061_),
    .Q(\_126_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13843_ (.CLK(clknet_leaf_94_clk),
    .D(_01062_),
    .Q(\_126_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13844_ (.CLK(clknet_leaf_93_clk),
    .D(_01063_),
    .Q(\_126_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13845_ (.CLK(clknet_leaf_93_clk),
    .D(_01064_),
    .Q(\_126_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13846_ (.CLK(clknet_leaf_92_clk),
    .D(_01065_),
    .Q(\_126_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13847_ (.CLK(clknet_leaf_92_clk),
    .D(_01066_),
    .Q(\_126_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13848_ (.CLK(clknet_leaf_90_clk),
    .D(_01067_),
    .Q(\_126_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13849_ (.CLK(clknet_leaf_90_clk),
    .D(_01068_),
    .Q(\_126_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13850_ (.CLK(clknet_leaf_89_clk),
    .D(_01069_),
    .Q(\_126_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13851_ (.CLK(clknet_leaf_72_clk),
    .D(_01070_),
    .Q(\_126_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13852_ (.CLK(clknet_leaf_71_clk),
    .D(_01071_),
    .Q(\_126_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13853_ (.CLK(clknet_leaf_72_clk),
    .D(_01072_),
    .Q(\_126_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13854_ (.CLK(clknet_leaf_69_clk),
    .D(_01073_),
    .Q(\_126_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13855_ (.CLK(clknet_leaf_65_clk),
    .D(_01074_),
    .Q(\_126_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13856_ (.CLK(clknet_leaf_64_clk),
    .D(_01075_),
    .Q(\_124_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13857_ (.CLK(clknet_leaf_69_clk),
    .D(_01076_),
    .Q(\_124_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13858_ (.CLK(clknet_leaf_65_clk),
    .D(_01077_),
    .Q(\_124_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13859_ (.CLK(clknet_leaf_64_clk),
    .D(_01078_),
    .Q(\_124_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13860_ (.CLK(clknet_leaf_63_clk),
    .D(_01079_),
    .Q(\_124_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13861_ (.CLK(clknet_leaf_64_clk),
    .D(_01080_),
    .Q(\_124_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13862_ (.CLK(clknet_leaf_62_clk),
    .D(_01081_),
    .Q(\_124_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13863_ (.CLK(clknet_leaf_62_clk),
    .D(_01082_),
    .Q(\_124_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13864_ (.CLK(clknet_leaf_62_clk),
    .D(_01083_),
    .Q(\_124_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13865_ (.CLK(clknet_leaf_62_clk),
    .D(_01084_),
    .Q(\_124_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13866_ (.CLK(clknet_leaf_97_clk),
    .D(_01085_),
    .Q(\_124_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13867_ (.CLK(clknet_leaf_95_clk),
    .D(_01086_),
    .Q(\_124_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13868_ (.CLK(clknet_leaf_97_clk),
    .D(_01087_),
    .Q(\_124_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13869_ (.CLK(clknet_leaf_97_clk),
    .D(_01088_),
    .Q(\_124_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13870_ (.CLK(clknet_leaf_98_clk),
    .D(_01089_),
    .Q(\_124_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13871_ (.CLK(clknet_leaf_95_clk),
    .D(_01090_),
    .Q(\_124_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13872_ (.CLK(clknet_leaf_96_clk),
    .D(_01091_),
    .Q(\_124_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13873_ (.CLK(clknet_leaf_95_clk),
    .D(_01092_),
    .Q(\_124_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13874_ (.CLK(clknet_leaf_96_clk),
    .D(_01093_),
    .Q(\_124_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13875_ (.CLK(clknet_leaf_95_clk),
    .D(_01094_),
    .Q(\_124_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13876_ (.CLK(clknet_leaf_92_clk),
    .D(_01095_),
    .Q(\_124_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13877_ (.CLK(clknet_leaf_93_clk),
    .D(_01096_),
    .Q(\_124_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13878_ (.CLK(clknet_leaf_92_clk),
    .D(_01097_),
    .Q(\_124_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13879_ (.CLK(clknet_leaf_92_clk),
    .D(_01098_),
    .Q(\_124_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13880_ (.CLK(clknet_leaf_90_clk),
    .D(_01099_),
    .Q(\_124_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13881_ (.CLK(clknet_leaf_90_clk),
    .D(_01100_),
    .Q(\_124_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13882_ (.CLK(clknet_leaf_89_clk),
    .D(_01101_),
    .Q(\_124_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13883_ (.CLK(clknet_leaf_89_clk),
    .D(_01102_),
    .Q(\_124_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13884_ (.CLK(clknet_leaf_72_clk),
    .D(_01103_),
    .Q(\_124_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13885_ (.CLK(clknet_leaf_72_clk),
    .D(_01104_),
    .Q(\_124_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13886_ (.CLK(clknet_leaf_69_clk),
    .D(_01105_),
    .Q(\_124_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13887_ (.CLK(clknet_leaf_69_clk),
    .D(_01106_),
    .Q(\_124_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13888_ (.CLK(clknet_leaf_69_clk),
    .D(_01107_),
    .Q(\_122_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13889_ (.CLK(clknet_leaf_69_clk),
    .D(_01108_),
    .Q(\_122_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13890_ (.CLK(clknet_leaf_64_clk),
    .D(_01109_),
    .Q(\_122_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13891_ (.CLK(clknet_leaf_64_clk),
    .D(_01110_),
    .Q(\_122_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13892_ (.CLK(clknet_leaf_64_clk),
    .D(_01111_),
    .Q(\_122_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13893_ (.CLK(clknet_leaf_64_clk),
    .D(_01112_),
    .Q(\_122_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13894_ (.CLK(clknet_leaf_64_clk),
    .D(_01113_),
    .Q(\_122_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13895_ (.CLK(clknet_leaf_64_clk),
    .D(_01114_),
    .Q(\_122_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13896_ (.CLK(clknet_leaf_64_clk),
    .D(_01115_),
    .Q(\_122_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13897_ (.CLK(clknet_leaf_64_clk),
    .D(_01116_),
    .Q(\_122_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13898_ (.CLK(clknet_leaf_97_clk),
    .D(_01117_),
    .Q(\_122_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13899_ (.CLK(clknet_leaf_95_clk),
    .D(_01118_),
    .Q(\_122_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13900_ (.CLK(clknet_leaf_97_clk),
    .D(_01119_),
    .Q(\_122_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13901_ (.CLK(clknet_leaf_97_clk),
    .D(_01120_),
    .Q(\_122_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13902_ (.CLK(clknet_leaf_98_clk),
    .D(_01121_),
    .Q(\_122_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13903_ (.CLK(clknet_leaf_97_clk),
    .D(_01122_),
    .Q(\_122_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13904_ (.CLK(clknet_leaf_96_clk),
    .D(_01123_),
    .Q(\_122_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13905_ (.CLK(clknet_leaf_95_clk),
    .D(_01124_),
    .Q(\_122_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13906_ (.CLK(clknet_leaf_96_clk),
    .D(_01125_),
    .Q(\_122_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13907_ (.CLK(clknet_leaf_95_clk),
    .D(_01126_),
    .Q(\_122_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13908_ (.CLK(clknet_leaf_92_clk),
    .D(_01127_),
    .Q(\_122_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13909_ (.CLK(clknet_leaf_93_clk),
    .D(_01128_),
    .Q(\_122_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13910_ (.CLK(clknet_leaf_96_clk),
    .D(_01129_),
    .Q(\_122_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13911_ (.CLK(clknet_leaf_92_clk),
    .D(_01130_),
    .Q(\_122_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13912_ (.CLK(clknet_leaf_91_clk),
    .D(_01131_),
    .Q(\_122_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13913_ (.CLK(clknet_leaf_91_clk),
    .D(_01132_),
    .Q(\_122_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13914_ (.CLK(clknet_leaf_91_clk),
    .D(_01133_),
    .Q(\_122_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13915_ (.CLK(clknet_leaf_90_clk),
    .D(_01134_),
    .Q(\_122_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13916_ (.CLK(clknet_leaf_72_clk),
    .D(_01135_),
    .Q(\_122_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13917_ (.CLK(clknet_leaf_72_clk),
    .D(_01136_),
    .Q(\_122_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13918_ (.CLK(clknet_leaf_68_clk),
    .D(_01137_),
    .Q(\_122_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13919_ (.CLK(clknet_leaf_69_clk),
    .D(_01138_),
    .Q(\_122_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13920_ (.CLK(clknet_leaf_70_clk),
    .D(_01139_),
    .Q(\_120_[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13921_ (.CLK(clknet_leaf_70_clk),
    .D(_01140_),
    .Q(\_120_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13922_ (.CLK(clknet_leaf_70_clk),
    .D(_01141_),
    .Q(\_120_[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13923_ (.CLK(clknet_leaf_70_clk),
    .D(_01142_),
    .Q(\_120_[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13924_ (.CLK(clknet_leaf_70_clk),
    .D(_01143_),
    .Q(\_120_[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13925_ (.CLK(clknet_leaf_70_clk),
    .D(_01144_),
    .Q(\_120_[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13926_ (.CLK(clknet_leaf_70_clk),
    .D(_01145_),
    .Q(\_120_[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13927_ (.CLK(clknet_leaf_70_clk),
    .D(_01146_),
    .Q(\_120_[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13928_ (.CLK(clknet_leaf_69_clk),
    .D(_01147_),
    .Q(\_120_[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13929_ (.CLK(clknet_leaf_69_clk),
    .D(_01148_),
    .Q(\_120_[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13930_ (.CLK(clknet_leaf_97_clk),
    .D(_01149_),
    .Q(\_120_[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13931_ (.CLK(clknet_leaf_96_clk),
    .D(_01150_),
    .Q(\_120_[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13932_ (.CLK(clknet_leaf_97_clk),
    .D(_01151_),
    .Q(\_120_[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13933_ (.CLK(clknet_leaf_97_clk),
    .D(_01152_),
    .Q(\_120_[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13934_ (.CLK(clknet_leaf_97_clk),
    .D(_01153_),
    .Q(\_120_[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13935_ (.CLK(clknet_leaf_97_clk),
    .D(_01154_),
    .Q(\_120_[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13936_ (.CLK(clknet_leaf_96_clk),
    .D(_01155_),
    .Q(\_120_[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13937_ (.CLK(clknet_leaf_95_clk),
    .D(_01156_),
    .Q(\_120_[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13938_ (.CLK(clknet_leaf_96_clk),
    .D(_01157_),
    .Q(\_120_[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13939_ (.CLK(clknet_leaf_96_clk),
    .D(_01158_),
    .Q(\_120_[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13940_ (.CLK(clknet_leaf_92_clk),
    .D(_01159_),
    .Q(\_120_[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13941_ (.CLK(clknet_leaf_93_clk),
    .D(_01160_),
    .Q(\_120_[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13942_ (.CLK(clknet_leaf_96_clk),
    .D(_01161_),
    .Q(\_120_[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13943_ (.CLK(clknet_leaf_91_clk),
    .D(_01162_),
    .Q(\_120_[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13944_ (.CLK(clknet_leaf_91_clk),
    .D(_01163_),
    .Q(\_120_[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13945_ (.CLK(clknet_leaf_91_clk),
    .D(_01164_),
    .Q(\_120_[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13946_ (.CLK(clknet_leaf_91_clk),
    .D(_01165_),
    .Q(\_120_[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13947_ (.CLK(clknet_leaf_90_clk),
    .D(_01166_),
    .Q(\_120_[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13948_ (.CLK(clknet_leaf_89_clk),
    .D(_01167_),
    .Q(\_120_[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13949_ (.CLK(clknet_leaf_90_clk),
    .D(_01168_),
    .Q(\_120_[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13950_ (.CLK(clknet_leaf_68_clk),
    .D(_01169_),
    .Q(\_120_[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13951_ (.CLK(clknet_leaf_69_clk),
    .D(_01170_),
    .Q(\_120_[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13952_ (.CLK(clknet_leaf_70_clk),
    .D(_01171_),
    .Q(\_118_[0] ));
 sky130_fd_sc_hd__dfxtp_2 _13953_ (.CLK(clknet_leaf_70_clk),
    .D(_01172_),
    .Q(\_118_[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13954_ (.CLK(clknet_leaf_71_clk),
    .D(_01173_),
    .Q(\_118_[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13955_ (.CLK(clknet_leaf_71_clk),
    .D(_01174_),
    .Q(\_118_[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13956_ (.CLK(clknet_leaf_71_clk),
    .D(_01175_),
    .Q(\_118_[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13957_ (.CLK(clknet_leaf_71_clk),
    .D(_01176_),
    .Q(\_118_[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13958_ (.CLK(clknet_leaf_72_clk),
    .D(_01177_),
    .Q(\_118_[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13959_ (.CLK(clknet_leaf_70_clk),
    .D(_01178_),
    .Q(\_118_[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13960_ (.CLK(clknet_leaf_71_clk),
    .D(_01179_),
    .Q(\_118_[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13961_ (.CLK(clknet_leaf_71_clk),
    .D(_01180_),
    .Q(\_118_[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13962_ (.CLK(clknet_leaf_97_clk),
    .D(_01181_),
    .Q(\_118_[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13963_ (.CLK(clknet_leaf_96_clk),
    .D(_01182_),
    .Q(\_118_[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13964_ (.CLK(clknet_leaf_97_clk),
    .D(_01183_),
    .Q(\_118_[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13965_ (.CLK(clknet_leaf_97_clk),
    .D(_01184_),
    .Q(\_118_[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13966_ (.CLK(clknet_leaf_97_clk),
    .D(_01185_),
    .Q(\_118_[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13967_ (.CLK(clknet_leaf_97_clk),
    .D(_01186_),
    .Q(\_118_[15] ));
 sky130_fd_sc_hd__dfxtp_4 _13968_ (.CLK(clknet_leaf_96_clk),
    .D(_01187_),
    .Q(\_118_[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13969_ (.CLK(clknet_leaf_96_clk),
    .D(_01188_),
    .Q(\_118_[17] ));
 sky130_fd_sc_hd__dfxtp_2 _13970_ (.CLK(clknet_leaf_96_clk),
    .D(_01189_),
    .Q(\_118_[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13971_ (.CLK(clknet_leaf_96_clk),
    .D(_01190_),
    .Q(\_118_[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13972_ (.CLK(clknet_leaf_93_clk),
    .D(_01191_),
    .Q(\_118_[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13973_ (.CLK(clknet_leaf_93_clk),
    .D(_01192_),
    .Q(\_118_[21] ));
 sky130_fd_sc_hd__dfxtp_2 _13974_ (.CLK(clknet_leaf_91_clk),
    .D(_01193_),
    .Q(\_118_[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13975_ (.CLK(clknet_leaf_92_clk),
    .D(_01194_),
    .Q(\_118_[23] ));
 sky130_fd_sc_hd__dfxtp_2 _13976_ (.CLK(clknet_leaf_91_clk),
    .D(_01195_),
    .Q(\_118_[24] ));
 sky130_fd_sc_hd__dfxtp_2 _13977_ (.CLK(clknet_leaf_91_clk),
    .D(_01196_),
    .Q(\_118_[25] ));
 sky130_fd_sc_hd__dfxtp_2 _13978_ (.CLK(clknet_leaf_91_clk),
    .D(_01197_),
    .Q(\_118_[26] ));
 sky130_fd_sc_hd__dfxtp_2 _13979_ (.CLK(clknet_leaf_90_clk),
    .D(_01198_),
    .Q(\_118_[27] ));
 sky130_fd_sc_hd__dfxtp_2 _13980_ (.CLK(clknet_leaf_90_clk),
    .D(_01199_),
    .Q(\_118_[28] ));
 sky130_fd_sc_hd__dfxtp_2 _13981_ (.CLK(clknet_leaf_90_clk),
    .D(_01200_),
    .Q(\_118_[29] ));
 sky130_fd_sc_hd__dfxtp_2 _13982_ (.CLK(clknet_leaf_68_clk),
    .D(_01201_),
    .Q(\_118_[30] ));
 sky130_fd_sc_hd__dfxtp_2 _13983_ (.CLK(clknet_leaf_68_clk),
    .D(_01202_),
    .Q(\_118_[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13984_ (.CLK(clknet_leaf_36_clk),
    .D(_01203_),
    .Q(_099_));
 sky130_fd_sc_hd__dfxtp_1 _13985_ (.CLK(clknet_leaf_31_clk),
    .D(_01204_),
    .Q(_096_));
 sky130_fd_sc_hd__dfxtp_1 _13986_ (.CLK(clknet_leaf_31_clk),
    .D(_01205_),
    .Q(_093_));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(din[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(din[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(din[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(din[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(din[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(din[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(din[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(din[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(din[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(din[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(din[19]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(din[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(din[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(din[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(din[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(din[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(din[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(din[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(din[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(din[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(din[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(din[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(din[2]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(din[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(din[31]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(din[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(din[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(din[5]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(din[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(din[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(din[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(din[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(dst_ready),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(rst),
    .X(net34));
 sky130_fd_sc_hd__buf_6 input35 (.A(src_ready),
    .X(net35));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(dout[0]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(dout[10]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(dout[11]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(dout[12]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(dout[13]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(dout[14]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(dout[15]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(dout[16]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(dout[17]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(dout[18]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(dout[19]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(dout[1]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(dout[20]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(dout[21]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(dout[22]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(dout[23]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(dout[24]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(dout[25]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(dout[26]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(dout[27]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(dout[28]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(dout[29]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(dout[2]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(dout[30]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(dout[31]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(dout[3]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(dout[4]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(dout[5]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(dout[6]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(dout[7]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(dout[8]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(dout[9]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(dst_write));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(src_read));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_1_0_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_1_0_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_1_1_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_1_1_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_opt_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_01274_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_01302_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_02353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_03667_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\_128_[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\_142_[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\_164_[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\_164_[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\_164_[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\_164_[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\_167_[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\_170_[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\_170_[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\_173_[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\_179_[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\_179_[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_01355_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_01519_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_01635_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_02001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_02001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_02237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_03568_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_04577_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(\_142_[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\_142_[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\_170_[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\_173_[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(\_173_[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\_179_[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\_182_[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(\_173_[7] ));
endmodule
