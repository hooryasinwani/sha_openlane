* NGSPICE file created from sha2_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt sha2_top VGND VPWR clk din[0] din[10] din[11] din[12] din[13] din[14] din[15]
+ din[16] din[17] din[18] din[19] din[1] din[20] din[21] din[22] din[23] din[24] din[25]
+ din[26] din[27] din[28] din[29] din[2] din[30] din[31] din[3] din[4] din[5] din[6]
+ din[7] din[8] din[9] dout[0] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15]
+ dout[16] dout[17] dout[18] dout[19] dout[1] dout[20] dout[21] dout[22] dout[23]
+ dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[2] dout[30] dout[31]
+ dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dst_ready dst_write rst
+ src_read src_ready
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09671_ _04049_ _04062_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__xor2_1
X_06883_ _243_\[29\] _01438_ _01513_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08622_ _02994_ _03021_ _03020_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__a21o_1
X_08553_ _185_\[3\] _02951_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__nand2_1
X_07504_ _182_\[12\] _01642_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__xor2_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08484_ _02890_ _02893_ _02916_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__o21a_1
XFILLER_35_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07435_ _01957_ _01987_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__or2_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07366_ _01918_ _01921_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__xnor2_4
XFILLER_108_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07297_ _01620_ _01827_ _01693_ _01855_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__a211o_1
X_09105_ _02262_ _03517_ _03518_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09036_ _02216_ _03418_ _03451_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__a21oi_1
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09938_ _04075_ _04005_ _04318_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__a21oi_1
XFILLER_104_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09869_ _03880_ _03927_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__nand2_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _118_\[31\] _120_\[31\] _01361_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__mux2_1
X_11900_ _152_\[16\] _05903_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__nand2_1
XFILLER_93_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11831_ _142_\[9\] _05841_ _05765_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__mux2_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11762_ _140_\[23\] _140_\[14\] VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__xnor2_1
X_13501_ clknet_leaf_36_clk _00720_ VGND VGND VPWR VPWR _158_\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _116_\[27\] _05704_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__nor2_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10713_ _167_\[11\] _04925_ _04938_ _04939_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__o211a_1
X_10644_ _176_\[22\] _04867_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__or2_1
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13432_ clknet_leaf_123_clk _00651_ VGND VGND VPWR VPWR _164_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10575_ _173_\[31\] _04836_ _04845_ _04839_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__a211o_1
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13363_ clknet_leaf_124_clk _00582_ VGND VGND VPWR VPWR _170_\[13\] sky130_fd_sc_hd__dfxtp_1
X_12314_ _06188_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13294_ clknet_leaf_26_clk _00513_ VGND VGND VPWR VPWR _176_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12245_ _06152_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__clkbuf_1
X_12176_ _06116_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11127_ _01258_ _05223_ _05194_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11058_ net51 _04628_ _05176_ _05117_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__o211a_1
X_10009_ _03893_ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__or2_1
XFILLER_76_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07220_ _01698_ _01780_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__xnor2_2
XFILLER_32_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07151_ _185_\[0\] _234_\[0\] VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__nand2_1
X_07082_ _237_\[17\] VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__clkbuf_8
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07984_ _02465_ _02499_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__nand2_1
X_09723_ _246_\[8\] _01314_ _03914_ _243_\[8\] _01455_ VGND VGND VPWR VPWR _04113_
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06935_ _240_\[11\] _01526_ _01510_ _01551_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__o211a_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09654_ _246_\[6\] _01313_ _01299_ _179_\[6\] VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__o22a_1
X_06866_ _243_\[24\] _01474_ _01461_ _01501_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__o211a_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08605_ _02830_ _02794_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__xnor2_1
X_09585_ _03901_ _03893_ _03979_ _03910_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__a211o_1
X_06797_ _01448_ _01450_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__or2_1
XFILLER_63_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08536_ _02964_ _02965_ _02967_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__o21a_1
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08467_ _228_\[1\] _231_\[1\] _02772_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__a21o_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07418_ _01965_ _01966_ _01971_ _01856_ _01884_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__a221oi_1
XFILLER_11_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08398_ net50 _02798_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__or2_1
X_07349_ _01904_ _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__nor2_2
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10360_ _04636_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__buf_4
XFILLER_136_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10291_ _182_\[7\] _04634_ _04647_ _04649_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__o211a_1
X_09019_ _03434_ _03435_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__nor2_1
X_12030_ _06010_ _06014_ _06008_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__o21ai_1
XFILLER_104_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13981_ clknet_leaf_90_clk _01200_ VGND VGND VPWR VPWR _118_\[29\] sky130_fd_sc_hd__dfxtp_2
X_12932_ clknet_leaf_39_clk _00151_ VGND VGND VPWR VPWR _246_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12863_ _06476_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _05804_ _05814_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__and2_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _06440_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__clkbuf_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _05760_ _05762_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__xnor2_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _149_\[26\] _05701_ _05625_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__mux2_1
X_13415_ clknet_leaf_12_clk _00634_ VGND VGND VPWR VPWR _164_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10627_ _02175_ _04818_ _04880_ _04823_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__o211a_1
XFILLER_127_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10558_ _01225_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__clkbuf_4
X_13346_ clknet_leaf_11_clk _00565_ VGND VGND VPWR VPWR _173_\[28\] sky130_fd_sc_hd__dfxtp_2
X_13277_ clknet_leaf_7_clk _00496_ VGND VGND VPWR VPWR _179_\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_142_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12228_ _06143_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__clkbuf_1
X_10489_ _01424_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__clkbuf_4
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12159_ _06107_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06720_ _01392_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06651_ _01351_ VGND VGND VPWR VPWR _436_\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_76_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06582_ _01289_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__clkbuf_1
X_09370_ _02862_ _01426_ _03379_ _03776_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__o211a_1
XFILLER_17_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08321_ _228_\[4\] _02771_ _02765_ _02783_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__o211a_1
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08252_ _01437_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07203_ _01752_ _01753_ _01763_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__or3_1
Xclkbuf_4_12_0_clk clknet_3_6_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_08183_ _234_\[30\] _02659_ _02636_ _02683_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__o211a_1
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07134_ _237_\[29\] VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__buf_6
X_07065_ _01645_ _01639_ _01609_ _01647_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__o211a_1
XFILLER_133_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07967_ _01856_ _02483_ _02502_ _02355_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__a211o_1
X_09706_ _04066_ _04069_ _04096_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__o21ai_1
X_06918_ _01448_ _01539_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__or2_1
XFILLER_74_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07898_ _02434_ _02435_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__nor2_1
X_09637_ _01235_ _03979_ _04026_ _04029_ _01230_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__o311a_1
X_06849_ _01448_ _01489_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__or2_1
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09568_ _195_\[5\] _03953_ _03956_ _03963_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__a31o_1
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08519_ _02852_ _02950_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__xnor2_2
X_09499_ _01282_ _03874_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__nor2b_4
XFILLER_130_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11530_ _05560_ _05562_ _05558_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11461_ _05508_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13200_ clknet_leaf_35_clk _00419_ VGND VGND VPWR VPWR _185_\[10\] sky130_fd_sc_hd__dfxtp_2
X_11392_ _05421_ _05428_ _05441_ _05445_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__and4bb_1
X_10412_ _179_\[16\] _04721_ _04705_ _04729_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__o211a_1
XFILLER_99_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10343_ _182_\[30\] _04678_ _04671_ _01710_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__a31o_1
X_13131_ clknet_leaf_117_clk _00350_ VGND VGND VPWR VPWR _228_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10274_ _179_\[1\] _04638_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__or2_1
X_13062_ clknet_leaf_112_clk _00281_ VGND VGND VPWR VPWR _234_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12013_ _140_\[11\] _140_\[13\] VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__xor2_1
XFILLER_78_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13964_ clknet_leaf_97_clk _01183_ VGND VGND VPWR VPWR _118_\[12\] sky130_fd_sc_hd__dfxtp_2
X_13895_ clknet_leaf_64_clk _01114_ VGND VGND VPWR VPWR _122_\[7\] sky130_fd_sc_hd__dfxtp_1
X_12915_ clknet_leaf_88_clk _00139_ VGND VGND VPWR VPWR _116_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12846_ _06467_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__clkbuf_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12777_ _06431_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__clkbuf_1
X_11728_ _05742_ _05745_ _05746_ _05747_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__a31o_1
XFILLER_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11659_ _118_\[28\] _118_\[0\] VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__xnor2_1
X_13329_ clknet_leaf_25_clk _00548_ VGND VGND VPWR VPWR _173_\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1_0_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_142_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08870_ _228_\[14\] _231_\[14\] _02814_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__a21o_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07821_ _01657_ _01608_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07752_ _01355_ _02282_ _02294_ _01884_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__a211o_1
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07683_ _182_\[17\] _01661_ _02169_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__a21o_1
X_06703_ _118_\[16\] _116_\[16\] _01381_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__mux2_1
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06634_ _01295_ _01252_ _01321_ _01332_ _01336_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__a2111o_1
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09422_ _228_\[30\] _231_\[30\] _02868_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__a21o_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09353_ _228_\[28\] _231_\[28\] _03759_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__o21a_1
X_06565_ _01273_ _01247_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__or2_4
XFILLER_80_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08304_ _228_\[0\] _02730_ _02753_ _02770_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__a211o_1
XFILLER_138_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06496_ _01207_ _01208_ _01209_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__or3_1
XFILLER_100_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09284_ _03630_ _03633_ _03692_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__a21o_1
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08235_ _164_\[13\] _02701_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__or2_1
XFILLER_121_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08166_ _02625_ _02671_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__or2_1
XFILLER_119_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07117_ _173_\[25\] _01646_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__or2_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08097_ _234_\[5\] _02564_ _02178_ _02622_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__a211o_1
XFILLER_133_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07048_ _240_\[9\] _01601_ _01598_ _01634_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__o211a_1
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08999_ _185_\[17\] _03383_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__nand2_1
XFILLER_56_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10961_ _164_\[20\] _167_\[20\] _01214_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__mux2_1
XFILLER_28_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12700_ _06391_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__clkbuf_1
X_13680_ clknet_leaf_78_clk _00899_ VGND VGND VPWR VPWR _136_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12631_ _126_\[8\] _124_\[8\] _06346_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__mux2_1
XFILLER_71_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10892_ _01424_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__clkbuf_4
XFILLER_12_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12562_ _128_\[7\] _126_\[7\] _06313_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__mux2_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12493_ _130_\[6\] _128_\[6\] _06280_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__mux2_1
X_11513_ _05555_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11444_ _118_\[10\] _118_\[6\] VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11375_ _149_\[26\] _132_\[26\] VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__nor2_1
XFILLER_140_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10326_ _182_\[23\] _04654_ _04642_ _04650_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__a31o_1
X_13114_ clknet_leaf_119_clk _00333_ VGND VGND VPWR VPWR _231_\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _03870_ _04622_ _04623_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13045_ clknet_leaf_108_clk _00264_ VGND VGND VPWR VPWR _237_\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10188_ _142_\[28\] _04557_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__and2_1
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13947_ clknet_leaf_90_clk _01166_ VGND VGND VPWR VPWR _120_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13878_ clknet_leaf_92_clk _01097_ VGND VGND VPWR VPWR _124_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12829_ _06458_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08020_ _02552_ _02553_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__nor2_1
XFILLER_128_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09971_ _04347_ _04350_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__nand2_1
XFILLER_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08922_ _185_\[15\] _03314_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__nand2_1
XFILLER_97_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08853_ _03272_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__xnor2_2
X_08784_ _03187_ _03188_ _03207_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__a21oi_1
X_07804_ _02281_ _02343_ _02344_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__a21bo_1
XFILLER_38_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07735_ _02277_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__inv_2
XFILLER_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07666_ _02209_ _02210_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__nand2_1
XFILLER_41_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09405_ _01519_ _03810_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__or2_1
XFILLER_37_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06617_ _01309_ _01311_ _01319_ _01295_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_111_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07597_ _02077_ _02102_ _02142_ _02143_ _02129_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__a311oi_4
XFILLER_41_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06548_ _158_\[7\] _158_\[8\] _01256_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__or3_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09336_ _02486_ _03714_ _03715_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__nand3_1
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09267_ _02862_ _03675_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__xnor2_1
X_08218_ _164_\[8\] _02701_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__or2_1
X_09198_ _03576_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__inv_2
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08149_ _167_\[20\] _231_\[20\] _02626_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__mux2_1
X_11160_ _01263_ _05248_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__nand2_1
XFILLER_136_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11091_ _158_\[0\] _05194_ _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__o21ai_1
XFILLER_121_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10111_ _142_\[23\] _04462_ _04463_ _04461_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__o2bb2ai_1
X_10042_ _03886_ _03983_ _04107_ _04418_ _01238_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__o311a_1
XFILLER_121_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13801_ clknet_leaf_60_clk _01020_ VGND VGND VPWR VPWR _128_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13732_ clknet_leaf_60_clk _00951_ VGND VGND VPWR VPWR _132_\[4\] sky130_fd_sc_hd__dfxtp_1
X_11993_ _05969_ _05987_ _05988_ _05950_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10944_ _167_\[15\] _05089_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__or2_1
X_13663_ clknet_leaf_55_clk _00882_ VGND VGND VPWR VPWR _138_\[31\] sky130_fd_sc_hd__dfxtp_1
X_10875_ _164_\[26\] _05025_ _05054_ _05035_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__a211o_1
XFILLER_31_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13594_ clknet_leaf_49_clk _00813_ VGND VGND VPWR VPWR _142_\[26\] sky130_fd_sc_hd__dfxtp_1
X_12614_ _01392_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12545_ _130_\[31\] _128_\[31\] _06302_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__mux2_1
XFILLER_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12476_ _132_\[30\] _130_\[30\] _06269_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__mux2_1
X_11427_ _149_\[0\] _05352_ _05477_ _05478_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__a22o_1
XANTENNA_5 _02359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11358_ _05416_ _05417_ _05409_ _05414_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__a211o_1
XFILLER_98_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10309_ _182_\[15\] _04654_ _04642_ _04650_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__a31o_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11289_ _152_\[14\] _05358_ _05318_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__mux2_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13028_ clknet_leaf_43_clk _00247_ VGND VGND VPWR VPWR _237_\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07520_ _02068_ _02069_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__nand2_1
XFILLER_47_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07451_ _01994_ _01995_ _02003_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__a21o_1
X_07382_ _01936_ _01937_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__or2_1
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09121_ _03499_ _03504_ _03497_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_123_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_123_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_129_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09052_ _170_\[20\] _02835_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__nor2_1
X_08003_ _01698_ _01827_ _02178_ _02537_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__a211o_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09954_ _04179_ _04215_ _04333_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__or3_1
X_09885_ _04268_ _04243_ _04244_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__o21ai_1
XFILLER_112_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08905_ _03323_ _03324_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__or2b_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08836_ _02071_ _03222_ _03257_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__o21a_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08767_ _02811_ _02772_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07718_ _01690_ _01645_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__xnor2_2
X_08698_ _03121_ _03124_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__xor2_1
XFILLER_26_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07649_ _02194_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__inv_2
X_10660_ _02535_ _04872_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__nand2_1
XFILLER_41_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09319_ _03724_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10591_ _04853_ _04854_ _04856_ _04839_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_114_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_114_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12330_ _136_\[25\] _134_\[25\] _06189_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__mux2_1
XFILLER_126_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12261_ _138_\[24\] _136_\[24\] _06156_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__mux2_1
XFILLER_107_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11212_ _152_\[4\] _05291_ _01362_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__mux2_1
XFILLER_107_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput42 net42 VGND VGND VPWR VPWR dout[15] sky130_fd_sc_hd__buf_2
X_12192_ _140_\[23\] _138_\[23\] _06123_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__mux2_1
Xoutput53 net53 VGND VGND VPWR VPWR dout[25] sky130_fd_sc_hd__buf_2
X_11143_ _05236_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__clkbuf_1
Xoutput64 net64 VGND VGND VPWR VPWR dout[6] sky130_fd_sc_hd__buf_2
XFILLER_1_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11074_ net57 _04848_ _05186_ _01436_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__a211o_1
X_10025_ _04399_ _04400_ _04396_ _04401_ _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__a221o_1
XFILLER_1_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11976_ _142_\[22\] _05262_ _05973_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__a21o_1
X_13715_ clknet_leaf_77_clk _00934_ VGND VGND VPWR VPWR _134_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10927_ net67 _05068_ _05091_ _05086_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__a211o_1
X_13646_ clknet_leaf_47_clk _00865_ VGND VGND VPWR VPWR _138_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10858_ _164_\[21\] _05025_ _05042_ _05035_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__a211o_1
X_13577_ clknet_leaf_52_clk _00796_ VGND VGND VPWR VPWR _142_\[9\] sky130_fd_sc_hd__dfxtp_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_105_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_105_clk sky130_fd_sc_hd__clkbuf_16
X_10789_ _167_\[2\] _170_\[2\] _04936_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__mux2_1
X_12528_ _130_\[23\] _128_\[23\] _06291_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__mux2_1
XFILLER_145_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12459_ _132_\[22\] _130_\[22\] _06258_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__mux2_1
XFILLER_113_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06951_ _176_\[16\] _01531_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__or2_1
X_09670_ _03871_ _04053_ _04054_ _04056_ _04061_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__a221o_1
XFILLER_95_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06882_ _179_\[29\] _01302_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__or2_1
XFILLER_82_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08621_ _03048_ _03049_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__xor2_2
XFILLER_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08552_ _01835_ _02982_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07503_ _02026_ _02027_ _02024_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__o21a_1
X_08483_ _185_\[1\] _02892_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__nand2_1
X_07434_ _01959_ _01960_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__and2b_1
XFILLER_62_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07365_ _01859_ _01862_ _01889_ _01920_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__o31a_2
XFILLER_10_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07296_ _01520_ _01833_ _01854_ _01799_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__o211a_1
X_09104_ _185_\[20\] _03484_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__and2_1
X_09035_ _03415_ _03417_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__nor2_1
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09937_ _01243_ _01284_ _03904_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__and3_1
XFILLER_77_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09868_ _04250_ _04251_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__nor2_1
XFILLER_85_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _04185_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__inv_2
XFILLER_93_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08819_ _03236_ _03240_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__or2_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11830_ _05839_ _05840_ net32 _05776_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11761_ _05770_ _05772_ _05769_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__a21o_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13500_ clknet_leaf_36_clk _00719_ VGND VGND VPWR VPWR _158_\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10712_ _01424_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__buf_2
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _05696_ _05707_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__or2_1
X_13431_ clknet_leaf_1_clk _00650_ VGND VGND VPWR VPWR _164_\[17\] sky130_fd_sc_hd__dfxtp_1
X_10643_ _02300_ _04818_ _04890_ _04891_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__o211a_1
X_10574_ _176_\[31\] _04833_ _04806_ _04844_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__o211a_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13362_ clknet_leaf_2_clk _00581_ VGND VGND VPWR VPWR _170_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12313_ _136_\[17\] _134_\[17\] _06178_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__mux2_1
XFILLER_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13293_ clknet_leaf_24_clk _00512_ VGND VGND VPWR VPWR _176_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12244_ _138_\[16\] _136_\[16\] _06145_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__mux2_1
XFILLER_123_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12175_ _140_\[15\] _138_\[15\] _06112_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__mux2_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11126_ _158_\[9\] _01257_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__nand2_1
XFILLER_95_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11057_ _04638_ _05175_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__or2_1
X_10008_ _04303_ _04385_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__nor2_1
XFILLER_45_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11959_ _140_\[31\] _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__xnor2_2
XFILLER_60_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13629_ clknet_leaf_51_clk _00848_ VGND VGND VPWR VPWR _140_\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07150_ _01687_ _01713_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__xnor2_2
X_07081_ _01421_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__buf_4
XFILLER_99_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09722_ _01231_ _04106_ _04109_ _04111_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__a211o_1
XFILLER_113_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07983_ _02516_ _02517_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__or2_1
X_06934_ _176_\[11\] _01531_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__or2_1
X_09653_ _243_\[6\] _03914_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__or2_1
X_06865_ _179_\[24\] _01301_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__or2_1
XFILLER_95_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09584_ _01241_ _03878_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__nor2_2
XFILLER_103_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08604_ _01867_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__inv_2
XFILLER_27_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06796_ _179_\[6\] _243_\[6\] _01449_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__mux2_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _02904_ _02928_ _02966_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__a21boi_1
XFILLER_36_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08466_ _02878_ _02899_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__xor2_1
XFILLER_51_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07417_ _01969_ _01970_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__xor2_4
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08397_ _225_\[22\] VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__buf_4
XFILLER_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07348_ _240_\[7\] _01626_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__and2b_1
XFILLER_124_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07279_ _01704_ _01837_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__xnor2_2
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10290_ _04648_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__clkbuf_4
X_09018_ _170_\[18\] _02827_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__and2_1
XFILLER_2_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13980_ clknet_leaf_90_clk _01199_ VGND VGND VPWR VPWR _118_\[28\] sky130_fd_sc_hd__dfxtp_2
XFILLER_58_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12931_ clknet_leaf_40_clk _00150_ VGND VGND VPWR VPWR _246_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12862_ _118_\[22\] _120_\[22\] _06473_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__mux2_1
XFILLER_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _05823_ _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__nand2_1
XFILLER_73_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _122_\[21\] _120_\[21\] _06434_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__mux2_1
XFILLER_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _05745_ _05752_ _05761_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__o21ai_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _05696_ _05700_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10626_ _04809_ _04879_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__or2_1
X_13414_ clknet_leaf_124_clk _00633_ VGND VGND VPWR VPWR _164_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13345_ clknet_leaf_10_clk _00564_ VGND VGND VPWR VPWR _173_\[27\] sky130_fd_sc_hd__dfxtp_2
X_10557_ _173_\[26\] _04818_ _04832_ _04823_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__o211a_1
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10488_ _04766_ _04783_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__or2_1
X_13276_ clknet_leaf_4_clk _00495_ VGND VGND VPWR VPWR _179_\[22\] sky130_fd_sc_hd__dfxtp_2
X_12227_ _138_\[8\] _136_\[8\] _06134_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__mux2_1
X_12158_ _140_\[7\] _138_\[7\] _06101_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__mux2_1
XFILLER_123_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12089_ _140_\[6\] _142_\[6\] _06068_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__mux2_1
X_11109_ _158_\[4\] _01254_ _158_\[5\] VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__o21ai_1
XFILLER_49_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06650_ _01327_ _01343_ _01341_ _01350_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__or4b_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06581_ _01287_ _01288_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__and2_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08320_ _02749_ _02782_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__or2_1
XFILLER_33_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08251_ _231_\[17\] _02730_ _02712_ _02732_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__a211o_1
XFILLER_20_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07202_ _01752_ _01753_ _01763_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08182_ _02625_ _02682_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__or2_1
XFILLER_118_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07133_ _240_\[28\] _01649_ _01693_ _01700_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__a211o_1
XFILLER_118_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07064_ _173_\[13\] _01646_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__or2_1
XFILLER_145_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07966_ _02500_ _02501_ _01354_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__o21a_1
X_09705_ _04063_ _04064_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__or2b_1
XFILLER_101_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06917_ _176_\[6\] _240_\[6\] _01449_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__mux2_1
XFILLER_55_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09636_ _03884_ _01292_ _04027_ _04028_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__o31ai_1
XFILLER_114_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07897_ _02389_ _02420_ _02432_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_94_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_16
X_06848_ _179_\[19\] _243_\[19\] _01449_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__mux2_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09567_ _03907_ _03959_ _03962_ _195_\[5\] VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__a211oi_1
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06779_ _01435_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__buf_4
X_09498_ _03891_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__clkbuf_4
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08518_ _02820_ _02784_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08449_ _170_\[0\] _02768_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__nand2_1
XFILLER_139_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11460_ _149_\[4\] _05507_ _05439_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__mux2_1
XFILLER_109_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11391_ _152_\[27\] _05262_ _05446_ _05447_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__a22o_1
X_10411_ _182_\[16\] _04696_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__or2_1
XFILLER_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10342_ _01217_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__buf_4
X_13130_ clknet_leaf_106_clk _00349_ VGND VGND VPWR VPWR _228_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13061_ clknet_leaf_110_clk _00280_ VGND VGND VPWR VPWR _234_\[5\] sky130_fd_sc_hd__dfxtp_1
X_12012_ _06006_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__clkbuf_1
X_10273_ _04637_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__buf_4
XFILLER_120_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_85_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13963_ clknet_leaf_96_clk _01182_ VGND VGND VPWR VPWR _118_\[11\] sky130_fd_sc_hd__dfxtp_2
X_13894_ clknet_leaf_64_clk _01113_ VGND VGND VPWR VPWR _122_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12914_ clknet_leaf_88_clk _00138_ VGND VGND VPWR VPWR _116_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12845_ _118_\[14\] _120_\[14\] _06462_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__mux2_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12776_ _122_\[13\] _120_\[13\] _06423_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__mux2_1
X_11727_ net1 _01274_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__and2_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11658_ _149_\[24\] _05352_ _05684_ _05685_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__a22o_1
XFILLER_127_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10609_ _02001_ _04868_ _04865_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__mux2_1
X_11589_ _05622_ _05623_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13328_ clknet_leaf_25_clk _00547_ VGND VGND VPWR VPWR _173_\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_143_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13259_ clknet_leaf_29_clk _00478_ VGND VGND VPWR VPWR _179_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07820_ _02336_ _02337_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__and2b_1
XFILLER_84_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07751_ _01778_ _02293_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_76_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_16
X_06702_ _01383_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__clkbuf_1
X_07682_ _02225_ _02226_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__nor2_2
XFILLER_53_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06633_ _01206_ _01329_ _01333_ _01328_ _01335_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__a221o_1
XFILLER_92_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09421_ _03788_ _03791_ _03824_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__nand3_1
X_06564_ _392_\[1\] _392_\[0\] VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__nor2_1
X_09352_ _228_\[28\] _231_\[28\] _02862_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__a21o_1
XFILLER_100_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08303_ _02768_ _02733_ _02760_ _02769_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__o211a_1
X_06495_ _392_\[4\] VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__inv_2
X_09283_ _03628_ _03659_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__nand2_1
X_08234_ _231_\[12\] _02690_ _02712_ _02720_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__a211o_1
X_08165_ _167_\[25\] _231_\[25\] _02626_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__mux2_1
XFILLER_134_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07116_ _237_\[25\] VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__buf_4
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08096_ _231_\[5\] _02611_ _01695_ _02621_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__o211a_1
XFILLER_134_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07047_ _01615_ _01633_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__or2_1
XFILLER_142_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08998_ _02249_ _03414_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_67_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07949_ _01623_ _01604_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__xnor2_2
XFILLER_56_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10960_ net46 _04853_ _05114_ _05067_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__o211a_1
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09619_ _04009_ _04012_ _03871_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__a21oi_1
X_10891_ _05028_ _05065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__or2_1
XFILLER_28_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12630_ _06354_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12561_ _06318_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__clkbuf_1
X_12492_ _06282_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__clkbuf_1
X_11512_ _149_\[9\] _05554_ _05533_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__mux2_1
XFILLER_8_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11443_ _05492_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11374_ _05432_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__clkbuf_1
X_13113_ clknet_leaf_103_clk _00332_ VGND VGND VPWR VPWR _231_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10325_ _179_\[22\] _04658_ _04668_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__a21o_1
X_10256_ _185_\[31\] _03868_ _03864_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__o21ai_1
X_13044_ clknet_leaf_108_clk _00263_ VGND VGND VPWR VPWR _237_\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10187_ _246_\[28\] _01316_ _04409_ _243_\[28\] _01511_ VGND VGND VPWR VPWR _04557_
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_58_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_120_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_11_0_clk clknet_3_5_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
X_13946_ clknet_leaf_91_clk _01165_ VGND VGND VPWR VPWR _120_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13877_ clknet_leaf_93_clk _01096_ VGND VGND VPWR VPWR _124_\[21\] sky130_fd_sc_hd__dfxtp_1
X_12828_ _118_\[6\] _120_\[6\] _06451_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__mux2_1
X_12759_ _122_\[5\] _120_\[5\] _06412_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__mux2_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09970_ _04308_ _04311_ _04348_ _04349_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__a31o_1
XFILLER_130_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08921_ _02817_ _03032_ _03309_ _03340_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__a211o_1
XFILLER_130_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08852_ _170_\[12\] _02807_ _03273_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__a21oi_1
XFILLER_97_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07803_ _02317_ _02313_ _02315_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_49_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_111_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08783_ _03205_ _03206_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__or2b_1
XFILLER_38_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07734_ _02195_ _02196_ _02276_ _02165_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__or4b_1
XFILLER_53_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07665_ _185_\[18\] _234_\[18\] VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__nand2_1
X_06616_ _093_ _01312_ _01317_ _01318_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__a211o_1
X_09404_ _03808_ _03809_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__xnor2_2
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07596_ _02132_ _02130_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__nor2_1
XFILLER_71_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06547_ _158_\[6\] _01255_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__or2_2
X_09335_ _02495_ _03720_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__nand2_1
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09266_ _02820_ _02790_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_opt_1_0_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_opt_1_0_clk sky130_fd_sc_hd__clkbuf_16
X_08217_ _231_\[7\] _02706_ _02695_ _02708_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__o211a_1
XFILLER_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09197_ _185_\[23\] _03575_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__nand2_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08148_ _01421_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__clkbuf_4
X_08079_ _01670_ _02609_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__or2_1
XFILLER_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11090_ _05195_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__buf_2
X_10110_ _04482_ _04483_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__nor2_1
X_10041_ _01243_ _01278_ _03873_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__or3b_1
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13800_ clknet_leaf_58_clk _01019_ VGND VGND VPWR VPWR _128_\[8\] sky130_fd_sc_hd__dfxtp_1
X_11992_ _05946_ _05961_ _05987_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__or3b_1
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13731_ clknet_leaf_60_clk _00950_ VGND VGND VPWR VPWR _132_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10943_ net41 _04853_ _05102_ _05067_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__o211a_1
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13662_ clknet_leaf_58_clk _00881_ VGND VGND VPWR VPWR _138_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10874_ _167_\[26\] _05022_ _05043_ _05053_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__o211a_1
Xclkbuf_3_0_0_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_13593_ clknet_leaf_49_clk _00812_ VGND VGND VPWR VPWR _142_\[25\] sky130_fd_sc_hd__dfxtp_1
X_12613_ _06345_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12544_ _06309_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12475_ _06273_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11426_ _116_\[0\] _05476_ _05263_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__o21a_1
XANTENNA_6 _02359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11357_ _05409_ _05414_ _05416_ _05417_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__o211a_1
XFILLER_125_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10308_ _179_\[14\] _04658_ _04659_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__a21o_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ clknet_leaf_17_clk _00246_ VGND VGND VPWR VPWR _237_\[3\] sky130_fd_sc_hd__dfxtp_1
X_11288_ _05356_ _05357_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__xnor2_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _04572_ _04568_ _04588_ _04589_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__o31a_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13929_ clknet_leaf_69_clk _01148_ VGND VGND VPWR VPWR _120_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07450_ _01923_ _02001_ _02002_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__a21o_1
XFILLER_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07381_ _01897_ _01928_ _01935_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__and3_1
XFILLER_50_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09120_ _03532_ _03533_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__and2_1
X_09051_ _02830_ _03032_ _03309_ _03466_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__a211o_1
XFILLER_129_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08002_ _02380_ _02526_ _02536_ _02202_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__o211a_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09953_ _03960_ _03907_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__nor2_1
XFILLER_103_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09884_ _04222_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__inv_2
XFILLER_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08904_ _03320_ _03322_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__nand2_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08835_ _185_\[12\] _03221_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__nand2_1
XFILLER_57_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08766_ _03167_ _03169_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__and2b_1
XFILLER_45_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07717_ _01667_ _01827_ _02178_ _02260_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__a211o_1
XFILLER_53_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08697_ _03122_ _03123_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__nand2_1
XFILLER_14_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07648_ _02158_ _02182_ _02193_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07579_ _243_\[15\] _240_\[15\] _01654_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__mux2_4
XFILLER_40_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09318_ _228_\[27\] _231_\[27\] _03725_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__o21a_1
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10590_ _01824_ _04855_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__nor2_1
XFILLER_126_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09249_ _03657_ _03658_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__and2_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12260_ _06160_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11211_ _05289_ _05290_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__xor2_1
X_12191_ _06124_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput43 net43 VGND VGND VPWR VPWR dout[16] sky130_fd_sc_hd__buf_2
XFILLER_135_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11142_ _05234_ _05235_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__or2_1
Xoutput54 net54 VGND VGND VPWR VPWR dout[26] sky130_fd_sc_hd__buf_2
Xoutput65 net65 VGND VGND VPWR VPWR dout[7] sky130_fd_sc_hd__buf_2
XFILLER_134_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11073_ _164_\[29\] _04872_ _04627_ _05185_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__o211a_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10024_ _04370_ _04371_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__and2b_1
XFILLER_102_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11975_ _05776_ _05971_ _05972_ _05263_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__o211a_1
XFILLER_91_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13714_ clknet_leaf_77_clk _00933_ VGND VGND VPWR VPWR _134_\[18\] sky130_fd_sc_hd__dfxtp_1
X_10926_ _164_\[9\] _05059_ _05043_ _05090_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__o211a_1
X_13645_ clknet_leaf_47_clk _00864_ VGND VGND VPWR VPWR _138_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10857_ _167_\[21\] _05022_ _05009_ _05041_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__o211a_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13576_ clknet_leaf_54_clk _00795_ VGND VGND VPWR VPWR _142_\[8\] sky130_fd_sc_hd__dfxtp_1
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10788_ _164_\[1\] _04986_ _04992_ _04952_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__a211o_1
XFILLER_9_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12527_ _06300_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__clkbuf_1
X_12458_ _06264_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11409_ _152_\[29\] _05279_ _05461_ _05463_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__o22a_1
XFILLER_141_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12389_ _06228_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06950_ _243_\[15\] _01536_ _01557_ _01562_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__a211o_1
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06881_ _246_\[28\] _01496_ _01509_ _01512_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__a211o_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08620_ _03015_ _03016_ _03017_ _03014_ _03012_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__o32ai_4
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08551_ _185_\[4\] _02981_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__xnor2_1
X_07502_ _02035_ _02052_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08482_ _02911_ _02914_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__xnor2_1
X_07433_ _01984_ _01985_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07364_ _182_\[7\] _01626_ _01919_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09103_ _185_\[20\] _03484_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__or2_1
X_07295_ _01852_ _01853_ _01427_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__a21o_1
X_09034_ _02252_ _03449_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09936_ _01237_ _04316_ _04253_ _01232_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__a31o_1
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09867_ _142_\[14\] _04249_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__nor2_1
XFILLER_97_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _01230_ _04178_ _04180_ _04182_ _04184_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__o32a_1
XFILLER_100_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08818_ _03236_ _03240_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__nand2_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08749_ _03136_ _03151_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__nand2_1
X_11760_ _01274_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__clkbuf_4
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10711_ _04888_ _04937_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__or2_1
XFILLER_26_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _05713_ _05714_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__nand2_1
XFILLER_14_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13430_ clknet_leaf_123_clk _00649_ VGND VGND VPWR VPWR _164_\[16\] sky130_fd_sc_hd__dfxtp_1
X_10642_ _01424_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10573_ _179_\[31\] _04799_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__or2_1
XFILLER_22_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13361_ clknet_leaf_0_clk _00580_ VGND VGND VPWR VPWR _170_\[11\] sky130_fd_sc_hd__dfxtp_1
X_13292_ clknet_leaf_26_clk _00511_ VGND VGND VPWR VPWR _176_\[6\] sky130_fd_sc_hd__dfxtp_1
X_12312_ _06187_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12243_ _06151_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12174_ _06115_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11125_ _158_\[8\] _05193_ _05221_ _05191_ _05222_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__a221o_1
XFILLER_49_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11056_ _164_\[23\] _03595_ _04636_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__mux2_1
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10007_ _03960_ _03952_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__nand2_1
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11958_ _140_\[6\] _140_\[8\] VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11889_ _05894_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__clkbuf_1
X_10909_ net62 _05048_ _05078_ _05067_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__o211a_1
X_13628_ clknet_leaf_51_clk _00847_ VGND VGND VPWR VPWR _140_\[28\] sky130_fd_sc_hd__dfxtp_2
XFILLER_60_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13559_ clknet_leaf_75_clk _00778_ VGND VGND VPWR VPWR _149_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07080_ _240_\[16\] _01649_ _01607_ _01659_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__a211o_1
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07982_ _02492_ _02504_ _02515_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__nor3_1
X_09721_ _01242_ _03897_ _04031_ _04110_ _04060_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__o311a_1
X_06933_ _243_\[10\] _01548_ _01545_ _01550_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__o211a_1
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09652_ _185_\[5\] _03869_ _03919_ _04044_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__o211a_1
XFILLER_103_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06864_ _246_\[23\] _01496_ _01460_ _01500_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__a211o_1
XFILLER_83_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09583_ _01235_ _03976_ _03977_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__nor3_1
X_06795_ _01339_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__buf_4
XFILLER_94_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08603_ _01406_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__clkbuf_4
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ _02925_ _02927_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__nand2_1
XFILLER_36_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08465_ _01734_ _02898_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__xnor2_1
X_07416_ _01918_ _01921_ _01917_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__o21ai_2
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08396_ _228_\[21\] _02838_ _02810_ _02841_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__a211o_1
XFILLER_137_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07347_ _01626_ _243_\[7\] VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__nor2_1
XFILLER_136_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07278_ _01657_ _01638_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__xnor2_1
X_09017_ _170_\[18\] _02827_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__nor2_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09919_ _03983_ _04138_ _04133_ _04300_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__o31a_1
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12930_ clknet_leaf_41_clk _00149_ VGND VGND VPWR VPWR _246_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12861_ _06475_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _152_\[8\] _05822_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__or2_1
XFILLER_73_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12792_ _06439_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__clkbuf_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _152_\[1\] _05751_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__nand2_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _05683_ _05697_ _05699_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__o21ai_1
XFILLER_42_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10625_ _173_\[16\] _176_\[16\] _04830_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__mux2_1
X_13413_ clknet_leaf_125_clk _00632_ VGND VGND VPWR VPWR _167_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10556_ _04809_ _04831_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__or2_1
X_13344_ clknet_leaf_12_clk _00563_ VGND VGND VPWR VPWR _173_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10487_ _176_\[6\] _179_\[6\] _04743_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__mux2_1
X_13275_ clknet_leaf_4_clk _00494_ VGND VGND VPWR VPWR _179_\[21\] sky130_fd_sc_hd__dfxtp_2
X_12226_ _06142_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12157_ _06106_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11108_ _05207_ _05208_ _05209_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__o21ai_1
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12088_ _06070_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11039_ _03376_ _04631_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__nor2_1
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06580_ _01239_ _01286_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__or2_1
XFILLER_80_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08250_ _228_\[17\] _02698_ _02723_ _02731_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__o211a_1
X_07201_ _01761_ _01762_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__xnor2_1
X_08181_ _167_\[30\] _231_\[30\] _02626_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__mux2_1
XFILLER_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07132_ _01698_ _01639_ _01695_ _01699_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__o211a_1
XFILLER_145_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07063_ _01339_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__clkbuf_2
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07965_ _02463_ _02470_ _02499_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__a21oi_1
X_09704_ _04093_ _04094_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__nand2_1
XFILLER_114_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06916_ _243_\[5\] _01536_ _01509_ _01538_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__a211o_1
X_09635_ _03884_ _04005_ _03933_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__a21oi_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07896_ _02433_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__inv_2
X_06847_ _246_\[18\] _01485_ _01481_ _01488_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__o211a_1
XFILLER_83_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09566_ _01240_ _03960_ _03961_ _01282_ _195_\[4\] VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__o221a_1
X_06778_ _01416_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__buf_4
XFILLER_71_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09497_ _03883_ _03887_ _03894_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__a21o_1
X_08517_ _01781_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__inv_2
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08448_ _02880_ _02882_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10410_ _176_\[15\] _04725_ _04727_ _04728_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__a211o_1
XFILLER_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08379_ net45 _02798_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__or2_1
XFILLER_137_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11390_ _05434_ _05442_ _05445_ _05263_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__o31a_1
XFILLER_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10341_ _182_\[29\] _04663_ _04676_ _04677_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__o211a_1
XFILLER_136_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13060_ clknet_leaf_110_clk _00279_ VGND VGND VPWR VPWR _234_\[4\] sky130_fd_sc_hd__dfxtp_1
X_10272_ _01214_ _04636_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__nor2_4
XFILLER_3_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12011_ _142_\[25\] _06003_ _06005_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__mux2_1
XFILLER_105_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13962_ clknet_leaf_97_clk _01181_ VGND VGND VPWR VPWR _118_\[10\] sky130_fd_sc_hd__dfxtp_2
X_12913_ clknet_leaf_88_clk _00137_ VGND VGND VPWR VPWR _116_\[22\] sky130_fd_sc_hd__dfxtp_1
X_13893_ clknet_leaf_64_clk _01112_ VGND VGND VPWR VPWR _122_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12844_ _06466_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12775_ _06430_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__clkbuf_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _152_\[0\] _05744_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__or2_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11657_ _05680_ _05683_ _05352_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10608_ _176_\[10\] _04867_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__or2_1
X_11588_ _05612_ _05614_ _05610_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__o21ai_1
XFILLER_115_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13327_ clknet_leaf_22_clk _00546_ VGND VGND VPWR VPWR _173_\[9\] sky130_fd_sc_hd__dfxtp_2
X_10539_ _04809_ _04819_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__or2_1
XFILLER_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13258_ clknet_leaf_29_clk _00477_ VGND VGND VPWR VPWR _179_\[4\] sky130_fd_sc_hd__dfxtp_1
X_13189_ clknet_leaf_33_clk _00408_ _00110_ VGND VGND VPWR VPWR _195_\[5\] sky130_fd_sc_hd__dfrtp_1
X_12209_ _06133_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07750_ _02291_ _02292_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__or2_2
X_06701_ _118_\[15\] _116_\[15\] _01381_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__mux2_1
XFILLER_80_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07681_ _182_\[18\] _01664_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__and2_1
X_06632_ _01207_ _01208_ _01334_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__and3b_1
XFILLER_53_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09420_ _03788_ _03791_ _03824_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__a21o_1
X_06563_ _392_\[4\] _01206_ _01251_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__or3_4
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09351_ _03756_ _03757_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__or2_1
X_09282_ _03689_ _03690_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__and2_1
X_08302_ net36 _02736_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__or2_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06494_ _392_\[3\] VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__buf_2
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08233_ _228_\[12\] _02698_ _02679_ _02719_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__o211a_1
XFILLER_21_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08164_ _234_\[24\] _02646_ _02664_ _02670_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__a211o_1
X_07115_ _240_\[24\] _01649_ _01607_ _01686_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__a211o_1
X_08095_ _167_\[5\] _02616_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__or2_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07046_ _173_\[9\] _01632_ _01617_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__mux2_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08997_ _185_\[18\] _03413_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__xnor2_1
X_07948_ _02459_ _02460_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__and2b_1
X_07879_ _02380_ _02403_ _02417_ _02202_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__o211a_1
X_09618_ _03952_ _04011_ _03872_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__o21ai_1
XFILLER_83_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10890_ _167_\[31\] _170_\[31\] _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__mux2_1
X_09549_ _03945_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__buf_2
XFILLER_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12560_ _128_\[6\] _126_\[6\] _06313_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__mux2_1
XFILLER_12_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12491_ _130_\[5\] _128_\[5\] _06280_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__mux2_1
X_11511_ _05552_ _05553_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__xnor2_1
X_11442_ _149_\[2\] _05491_ _05439_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__mux2_1
XFILLER_109_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11373_ _152_\[25\] _05431_ _05318_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__mux2_1
XFILLER_124_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10324_ _182_\[22\] _04654_ _04642_ _04650_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__a31o_1
X_13112_ clknet_leaf_103_clk _00331_ VGND VGND VPWR VPWR _231_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10255_ _04610_ _04621_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13043_ clknet_leaf_110_clk _00262_ VGND VGND VPWR VPWR _237_\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10186_ _04533_ _04555_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__and2_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13945_ clknet_leaf_91_clk _01164_ VGND VGND VPWR VPWR _120_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13876_ clknet_leaf_92_clk _01095_ VGND VGND VPWR VPWR _124_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12827_ _06457_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12758_ _06421_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__clkbuf_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12689_ _06385_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__clkbuf_1
X_11709_ _05715_ _05719_ _05726_ _05713_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__o211ai_2
XFILLER_30_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08920_ _01409_ _03332_ _03333_ _03339_ _01799_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__o311a_1
XFILLER_123_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08851_ _03210_ _03246_ _03245_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__o21ba_1
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07802_ _02342_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__inv_2
X_08782_ _03189_ _03190_ _03204_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__o21ai_1
X_07733_ _02220_ _02256_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__nand2_1
XFILLER_38_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07664_ _185_\[18\] _234_\[18\] VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__or2_1
XFILLER_38_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06615_ _01206_ _01247_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__nor2_2
XFILLER_111_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09403_ _03770_ _03771_ _03772_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__a21bo_1
XFILLER_25_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07595_ _02101_ _02131_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__and2_1
X_06546_ _158_\[5\] _158_\[4\] _01254_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__or3_1
XFILLER_40_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09334_ _03724_ _03726_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__and2b_1
XFILLER_139_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09265_ _02422_ _03673_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__nand2_1
X_09196_ _03600_ _03606_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__xor2_2
X_08216_ _02686_ _02707_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__or2_1
XFILLER_119_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08147_ _234_\[19\] _02646_ _02629_ _02658_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__a211o_1
XFILLER_134_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08078_ _167_\[0\] _231_\[0\] _01672_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__mux2_1
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07029_ _237_\[5\] VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__buf_4
X_10040_ _04280_ _04416_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__or2_1
XFILLER_103_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11991_ _05968_ _05978_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__nor2_1
XFILLER_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13730_ clknet_leaf_59_clk _00949_ VGND VGND VPWR VPWR _132_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10942_ _05079_ _05101_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__or2_1
XFILLER_29_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13661_ clknet_leaf_56_clk _00880_ VGND VGND VPWR VPWR _138_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10873_ _170_\[26\] _05036_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__or2_1
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12612_ _128_\[31\] _126_\[31\] _06335_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__mux2_1
X_13592_ clknet_leaf_50_clk _00811_ VGND VGND VPWR VPWR _142_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12543_ _130_\[30\] _128_\[30\] _06302_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__mux2_1
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12474_ _132_\[29\] _130_\[29\] _06269_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__mux2_1
X_11425_ _116_\[0\] _05476_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__nand2_1
XANTENNA_7 _02416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11356_ _149_\[23\] _132_\[23\] VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__nand2_1
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10307_ _182_\[14\] _04654_ _04642_ _04650_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__a31o_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13026_ clknet_leaf_17_clk _00245_ VGND VGND VPWR VPWR _237_\[2\] sky130_fd_sc_hd__dfxtp_1
X_11287_ _05342_ _05344_ _05349_ _05348_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__a31o_1
XFILLER_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10238_ _04604_ _04605_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__and2b_1
XFILLER_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10169_ _04103_ _03878_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__nor2_1
XFILLER_67_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13928_ clknet_leaf_69_clk _01147_ VGND VGND VPWR VPWR _120_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13859_ clknet_leaf_64_clk _01078_ VGND VGND VPWR VPWR _124_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07380_ _01897_ _01928_ _01935_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__a21oi_1
X_09050_ _01409_ _03460_ _03461_ _03465_ _01799_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__o311a_1
XFILLER_129_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08001_ _02404_ _02535_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__nand2_1
XFILLER_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09952_ _185_\[17\] _04150_ _04175_ _04332_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__o211a_1
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08903_ _03320_ _03322_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__nor2_1
X_09883_ _04224_ _04243_ _04244_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__or3b_1
XFILLER_112_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08834_ _02064_ _03255_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08765_ _03164_ _03166_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__nor2_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07716_ _01520_ _02237_ _02259_ _02202_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__o211a_1
XFILLER_38_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08696_ _03025_ _03054_ _03058_ _03064_ _03066_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__a311o_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07647_ _02191_ _02192_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07578_ _02123_ _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06529_ _01237_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__buf_2
X_09317_ _228_\[27\] _231_\[27\] _02858_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__a21o_1
XFILLER_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09248_ _03638_ _03639_ _03656_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__or3_1
XFILLER_31_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09179_ _03589_ _03590_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_10_0_clk clknet_3_5_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
X_11210_ _05274_ _05280_ _05283_ _05281_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__o31a_1
X_12190_ _140_\[22\] _138_\[22\] _06123_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__mux2_1
XFILLER_31_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11141_ net14 _05190_ _05192_ _158_\[12\] VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__a22o_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput66 net66 VGND VGND VPWR VPWR dout[8] sky130_fd_sc_hd__buf_2
Xoutput44 net44 VGND VGND VPWR VPWR dout[17] sky130_fd_sc_hd__buf_2
Xoutput55 net55 VGND VGND VPWR VPWR dout[27] sky130_fd_sc_hd__buf_2
X_11072_ _03810_ _04625_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__or2_1
XFILLER_0_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10023_ _04308_ _04348_ _04349_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11974_ net15 _05742_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__or2_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13713_ clknet_leaf_77_clk _00932_ VGND VGND VPWR VPWR _134_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10925_ _167_\[9\] _05089_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__or2_1
XFILLER_112_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13644_ clknet_leaf_78_clk _00863_ VGND VGND VPWR VPWR _138_\[12\] sky130_fd_sc_hd__dfxtp_1
X_10856_ _170_\[21\] _05036_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__or2_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13575_ clknet_leaf_54_clk _00794_ VGND VGND VPWR VPWR _142_\[7\] sky130_fd_sc_hd__dfxtp_2
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10787_ _167_\[1\] _04980_ _04958_ _04991_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__o211a_1
XFILLER_40_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12526_ _130_\[22\] _128_\[22\] _06291_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__mux2_1
X_12457_ _132_\[21\] _130_\[21\] _06258_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__mux2_1
XFILLER_8_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11408_ _05263_ _05462_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__nand2_1
XFILLER_126_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12388_ _132_\[20\] _134_\[20\] _06219_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__mux2_1
XFILLER_140_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11339_ _149_\[21\] _132_\[21\] VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__nor2_1
XFILLER_141_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06880_ _243_\[28\] _01474_ _01510_ _01511_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__o211a_1
XFILLER_79_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13009_ clknet_leaf_10_clk _00228_ VGND VGND VPWR VPWR _240_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08550_ _02855_ _02980_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__xnor2_2
X_07501_ _02050_ _02051_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__nor2_1
X_08481_ _185_\[2\] _02913_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07432_ _243_\[10\] _240_\[10\] _01635_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__mux2_2
XFILLER_63_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07363_ _182_\[6\] _01623_ _01887_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__and3_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09102_ _03514_ _03515_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__nand2_1
X_07294_ _01849_ _01850_ _01851_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__or3_1
XFILLER_108_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09033_ _03446_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09935_ _04075_ _03890_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__nand2_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09866_ _142_\[14\] _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__and2_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08817_ _03100_ _03238_ _03239_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__o21ai_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _03872_ _04183_ _01230_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__o21ai_1
XFILLER_100_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08748_ _03117_ _03152_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__nand2_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _185_\[7\] _03072_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__nand2_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10710_ _170_\[11\] _173_\[11\] _04936_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__mux2_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _116_\[28\] _05712_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__or2_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10641_ _04888_ _04889_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__or2_1
X_10572_ _173_\[30\] _04818_ _04843_ _04823_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__o211a_1
X_13360_ clknet_leaf_2_clk _00579_ VGND VGND VPWR VPWR _170_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12311_ _136_\[16\] _134_\[16\] _06178_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__mux2_1
X_13291_ clknet_leaf_26_clk _00510_ VGND VGND VPWR VPWR _176_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12242_ _138_\[15\] _136_\[15\] _06145_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__mux2_1
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12173_ _140_\[14\] _138_\[14\] _06112_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__mux2_1
XFILLER_123_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11124_ net9 _05190_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__and2_1
XFILLER_96_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11055_ _03544_ _04861_ _05174_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__a21boi_1
X_10006_ _01244_ _01281_ _04383_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__a21o_1
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11957_ _05944_ _05955_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__nand2_1
XFILLER_45_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10908_ _05028_ _05077_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__or2_1
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11888_ _142_\[14\] _05892_ _05893_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__mux2_1
XFILLER_60_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13627_ clknet_leaf_50_clk _00846_ VGND VGND VPWR VPWR _140_\[27\] sky130_fd_sc_hd__dfxtp_2
XFILLER_60_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10839_ _167_\[16\] _170_\[16\] _04995_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__mux2_1
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13558_ clknet_leaf_76_clk _00777_ VGND VGND VPWR VPWR _149_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12509_ _06200_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__clkbuf_4
XFILLER_9_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13489_ clknet_leaf_42_clk _00708_ VGND VGND VPWR VPWR _158_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07981_ _02492_ _02504_ _02515_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__o21a_1
X_09720_ _04081_ _04010_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__or2_1
XFILLER_113_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06932_ _01448_ _01549_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__or2_1
XFILLER_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09651_ _04042_ _04043_ _03868_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06863_ _243_\[23\] _01474_ _01461_ _01499_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__o211a_1
XFILLER_83_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09582_ _01241_ _03888_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__nand2_1
XFILLER_103_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06794_ _01405_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__buf_2
X_08602_ _02784_ _02838_ _02861_ _03031_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__a211o_1
XFILLER_82_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08533_ _02947_ _02948_ _02963_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__nor3_1
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08464_ _02894_ _02897_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__xor2_1
X_07415_ _01967_ _01968_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__nand2_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08395_ _02839_ _02791_ _02824_ _02840_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__o211a_1
X_07346_ _01901_ _01902_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__or2_1
XFILLER_109_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07277_ _01835_ _01809_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__or2_1
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09016_ _03428_ _03431_ _01523_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__o21a_1
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09918_ _03880_ _03984_ _04132_ _01237_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__a211o_1
XFILLER_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09849_ _03871_ _03925_ _04233_ _04078_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__a31o_1
XFILLER_100_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12860_ _118_\[21\] _120_\[21\] _06473_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__mux2_1
XFILLER_37_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _152_\[8\] _05822_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__nand2_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12791_ _122_\[20\] _120_\[20\] _06434_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__mux2_1
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _05758_ _05759_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__nand2_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _116_\[25\] _05687_ _05698_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__a21oi_1
XFILLER_139_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10624_ _02139_ _04861_ _04878_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__a21boi_1
X_13412_ clknet_leaf_128_clk _00631_ VGND VGND VPWR VPWR _167_\[30\] sky130_fd_sc_hd__dfxtp_2
X_13343_ clknet_leaf_11_clk _00562_ VGND VGND VPWR VPWR _173_\[25\] sky130_fd_sc_hd__dfxtp_2
X_10555_ _176_\[26\] _179_\[26\] _04830_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__mux2_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10486_ _173_\[5\] _04780_ _04782_ _04740_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__o211a_1
XFILLER_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13274_ clknet_leaf_4_clk _00493_ VGND VGND VPWR VPWR _179_\[20\] sky130_fd_sc_hd__dfxtp_2
X_12225_ _138_\[7\] _136_\[7\] _06134_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__mux2_1
XFILLER_108_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12156_ _140_\[6\] _138_\[6\] _06101_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__mux2_1
X_11107_ _01254_ _05194_ _05196_ _158_\[4\] VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__o211ai_1
XFILLER_110_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12087_ _140_\[5\] _142_\[5\] _06068_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__mux2_1
XFILLER_110_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11038_ net43 _164_\[16\] _01215_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__mux2_1
XFILLER_64_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12989_ clknet_leaf_22_clk _00208_ VGND VGND VPWR VPWR _243_\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_45_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07200_ _243_\[2\] _240_\[2\] _01608_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__mux2_2
X_08180_ _234_\[29\] _02646_ _02664_ _02681_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__a211o_1
XFILLER_32_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07131_ _173_\[28\] _01646_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__or2_1
XFILLER_145_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07062_ _237_\[13\] VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__buf_6
XFILLER_114_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07964_ _02463_ _02470_ _02499_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__and3_1
X_09703_ _04047_ _04072_ _04092_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__or3_1
X_06915_ _240_\[5\] _01526_ _01510_ _01537_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__o211a_1
XFILLER_56_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07895_ _02389_ _02420_ _02432_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__o21ai_1
X_09634_ _01280_ _03888_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__nor2_1
X_06846_ _01444_ _01487_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__nand2_1
XFILLER_83_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09565_ _01277_ _01279_ _195_\[3\] VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__o21ba_1
X_06777_ _246_\[2\] _01422_ _01425_ _01434_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__o211a_1
XFILLER_71_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09496_ _03888_ _03893_ _01234_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__a21o_1
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08516_ _02922_ _02924_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__and2b_1
XFILLER_23_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08447_ _228_\[0\] _231_\[0\] _02881_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__o21a_1
XFILLER_11_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08378_ _225_\[18\] VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__buf_4
X_07329_ _01480_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__buf_4
XFILLER_109_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10340_ _01424_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10271_ _04635_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__buf_4
X_12010_ _06004_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__buf_4
XFILLER_3_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13961_ clknet_leaf_71_clk _01180_ VGND VGND VPWR VPWR _118_\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12912_ clknet_leaf_88_clk _00136_ VGND VGND VPWR VPWR _116_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13892_ clknet_leaf_64_clk _01111_ VGND VGND VPWR VPWR _122_\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12843_ _118_\[13\] _120_\[13\] _06462_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__mux2_1
XFILLER_27_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12774_ _122_\[12\] _120_\[12\] _06423_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__mux2_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _152_\[0\] _05744_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__nand2_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11656_ _05680_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__or2_1
XFILLER_30_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10607_ _01212_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__buf_4
X_11587_ _05619_ _05621_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__nand2_1
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13326_ clknet_leaf_25_clk _00545_ VGND VGND VPWR VPWR _173_\[8\] sky130_fd_sc_hd__dfxtp_2
X_10538_ _176_\[21\] _179_\[21\] _04790_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__mux2_1
X_13257_ clknet_leaf_24_clk _00476_ VGND VGND VPWR VPWR _179_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12208_ _140_\[31\] _138_\[31\] _06123_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__mux2_1
X_10469_ _04766_ _04769_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__or2_1
X_13188_ clknet_leaf_33_clk _00407_ _00109_ VGND VGND VPWR VPWR _195_\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12139_ _140_\[30\] _142_\[30\] _06090_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__mux2_1
XFILLER_111_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06700_ _01382_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07680_ _182_\[18\] _01664_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__nor2_1
X_06631_ _096_ _01306_ _01268_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06562_ _01266_ _01270_ _01249_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__a21oi_2
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09350_ _03718_ _03742_ _03755_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__and3_1
X_09281_ _03651_ _03670_ _03688_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__or3_1
XFILLER_21_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08301_ _225_\[0\] VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__buf_4
X_06493_ _392_\[2\] VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__buf_2
XFILLER_21_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08232_ _164_\[12\] _02701_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__or2_1
XFILLER_119_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08163_ _231_\[24\] _02649_ _02641_ _02669_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__o211a_1
XFILLER_119_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07114_ _01684_ _01639_ _01609_ _01685_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__o211a_1
X_08094_ _234_\[4\] _02564_ _02178_ _02620_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__a211o_1
XFILLER_9_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07045_ _237_\[9\] VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__buf_6
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08996_ _02871_ _03412_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__xnor2_2
XFILLER_125_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07947_ _02481_ _02482_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__xor2_2
X_07878_ _02404_ _02416_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__nand2_1
XFILLER_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09617_ _04010_ _03977_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__nor2_1
X_06829_ _01427_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__clkbuf_4
XFILLER_71_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09548_ _01275_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__clkbuf_4
XFILLER_55_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09479_ _195_\[1\] _195_\[0\] VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__xor2_1
X_11510_ _05539_ _05544_ _05542_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12490_ _06281_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11441_ _05488_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11372_ _05428_ _05430_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10323_ _179_\[21\] _04658_ _04667_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__a21o_1
X_13111_ clknet_leaf_103_clk _00330_ VGND VGND VPWR VPWR _231_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10254_ _04612_ _04620_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13042_ clknet_leaf_110_clk _00261_ VGND VGND VPWR VPWR _237_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10185_ _04527_ _04548_ _04549_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__o21ba_1
XFILLER_105_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13944_ clknet_leaf_91_clk _01163_ VGND VGND VPWR VPWR _120_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13875_ clknet_leaf_95_clk _01094_ VGND VGND VPWR VPWR _124_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12826_ _118_\[5\] _120_\[5\] _06451_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__mux2_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12757_ _122_\[4\] _120_\[4\] _06412_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__mux2_1
XFILLER_91_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12688_ _124_\[3\] _122_\[3\] _06379_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__mux2_1
X_11708_ _05730_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__clkbuf_1
X_11639_ _149_\[22\] _05668_ _05625_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__mux2_1
XFILLER_30_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13309_ clknet_leaf_4_clk _00528_ VGND VGND VPWR VPWR _176_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08850_ _03270_ _03271_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__nand2_1
XFILLER_111_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07801_ _02275_ _02316_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__nand2_1
X_08781_ _03189_ _03190_ _03204_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__nor3_1
XFILLER_84_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07732_ _02272_ _02274_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__xnor2_1
X_07663_ _01701_ _02207_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__xnor2_2
XFILLER_38_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06614_ _01316_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__inv_2
XFILLER_111_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09402_ _03806_ _03807_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__nand2_1
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07594_ _01654_ _01973_ _01886_ _02141_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__o211a_1
X_09333_ _03630_ _03633_ _03692_ _03738_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__a211o_1
XFILLER_25_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06545_ _158_\[1\] _158_\[0\] _158_\[3\] _158_\[2\] VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_126_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_126_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09264_ _03645_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__inv_2
XFILLER_138_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09195_ _03375_ _03470_ _03601_ _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__o31a_1
X_08215_ _164_\[7\] _228_\[7\] _02687_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__mux2_1
X_08146_ _231_\[19\] _02649_ _02641_ _02657_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__o211a_1
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08077_ _01707_ _02448_ _02419_ _02608_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__o211a_1
XFILLER_106_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07028_ _240_\[4\] _01601_ _01598_ _01619_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__o211a_1
XFILLER_121_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08979_ _03396_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__inv_2
XFILLER_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11990_ _05984_ _05985_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__nand2_1
XFILLER_91_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10941_ _164_\[14\] _167_\[14\] _05064_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__mux2_1
X_13660_ clknet_leaf_56_clk _00879_ VGND VGND VPWR VPWR _138_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12611_ _06344_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10872_ _164_\[25\] _05048_ _05052_ _04998_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__o211a_1
X_13591_ clknet_leaf_46_clk _00810_ VGND VGND VPWR VPWR _142_\[23\] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_117_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_117_clk sky130_fd_sc_hd__clkbuf_16
X_12542_ _06308_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12473_ _06272_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11424_ _118_\[18\] _05475_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_8 _02645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11355_ _149_\[23\] _132_\[23\] VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__or2_1
X_11286_ _05354_ _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__and2_1
X_10306_ _04633_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__clkbuf_4
X_10237_ _04582_ _04585_ _04603_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__or3b_1
X_13025_ clknet_leaf_17_clk _00244_ VGND VGND VPWR VPWR _237_\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10168_ _142_\[27\] _04538_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10099_ _142_\[24\] _04471_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__nor2_1
X_13927_ clknet_leaf_70_clk _01146_ VGND VGND VPWR VPWR _120_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13858_ clknet_leaf_65_clk _01077_ VGND VGND VPWR VPWR _124_\[2\] sky130_fd_sc_hd__dfxtp_1
X_13789_ clknet_leaf_69_clk _01008_ VGND VGND VPWR VPWR _130_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12809_ _122_\[29\] _120_\[29\] _01367_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_108_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_108_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_43_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08000_ _02531_ _02534_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__xnor2_2
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09951_ _03945_ _04330_ _04331_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__or3_1
XFILLER_143_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08902_ _02097_ _03284_ _03321_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__a21oi_1
X_09882_ _04264_ _04265_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08833_ _185_\[13\] _03254_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08764_ _03172_ _03177_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__nand2_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07715_ _02257_ _02258_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__or2_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08695_ _170_\[7\] _02790_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__or2_1
XFILLER_26_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07646_ _243_\[17\] _240_\[17\] _01661_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__mux2_4
XFILLER_53_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07577_ _02124_ _02092_ _02091_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__o21a_1
XFILLER_13_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06528_ _01236_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__buf_2
X_09316_ _03722_ _03723_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__or2_1
X_09247_ _03638_ _03639_ _03656_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__o21ai_1
XFILLER_31_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09178_ _03564_ _03567_ _03562_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__a21bo_1
X_08129_ _234_\[14\] _02564_ _02629_ _02645_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__a211o_1
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11140_ _01260_ _05233_ _05194_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__a21oi_1
Xoutput67 net67 VGND VGND VPWR VPWR dout[9] sky130_fd_sc_hd__buf_2
XFILLER_134_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput56 net56 VGND VGND VPWR VPWR dout[28] sky130_fd_sc_hd__buf_2
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput45 net45 VGND VGND VPWR VPWR dout[18] sky130_fd_sc_hd__buf_2
XFILLER_89_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11071_ net56 _04628_ _05184_ _05117_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__o211a_1
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10022_ _04371_ _04370_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__or2b_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11973_ _05968_ _05970_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13712_ clknet_leaf_78_clk _00931_ VGND VGND VPWR VPWR _134_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10924_ _01216_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__clkbuf_2
X_13643_ clknet_leaf_48_clk _00862_ VGND VGND VPWR VPWR _138_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10855_ _164_\[20\] _04983_ _05040_ _04998_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__o211a_1
X_13574_ clknet_leaf_34_clk _00793_ VGND VGND VPWR VPWR _142_\[6\] sky130_fd_sc_hd__dfxtp_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _06299_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10786_ _170_\[1\] _04953_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__or2_1
XFILLER_12_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12456_ _06263_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11407_ _05458_ _05459_ _05460_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__a21o_1
X_12387_ _06227_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11338_ _05279_ _05399_ _05400_ _05401_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__a31o_1
XFILLER_140_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11269_ _149_\[12\] _132_\[12\] VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__or2_1
XFILLER_100_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13008_ clknet_leaf_14_clk _00227_ VGND VGND VPWR VPWR _240_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07500_ _02014_ _02036_ _02049_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__nor3_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08480_ _02849_ _02912_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__xnor2_1
X_07431_ _01982_ _01983_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__nand2_1
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07362_ _01916_ _01917_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__nand2_2
XFILLER_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09101_ _02271_ _03489_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__nand2_1
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07293_ _01849_ _01850_ _01851_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__o21ai_1
XFILLER_31_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09032_ _02249_ _03414_ _03447_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__o21ai_1
XFILLER_129_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09934_ _01237_ _04314_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__nor2_1
XFILLER_89_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09865_ _246_\[14\] _01314_ _04129_ _243_\[14\] _01472_ VGND VGND VPWR VPWR _04249_
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08816_ _03187_ _03205_ _03237_ _03176_ _03206_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__o221a_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _04055_ _04080_ _03928_ _03880_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__a22o_1
XFILLER_133_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08747_ _03170_ _03171_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__xor2_1
XFILLER_39_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _03101_ _03104_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__xnor2_4
XFILLER_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _01923_ _02175_ _02002_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__a21o_1
XFILLER_54_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10640_ _173_\[21\] _176_\[21\] _04830_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__mux2_1
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10571_ _04809_ _04842_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__or2_1
X_12310_ _06186_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__clkbuf_1
X_13290_ clknet_leaf_24_clk _00509_ VGND VGND VPWR VPWR _176_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12241_ _06150_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12172_ _06114_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11123_ _01257_ _05220_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__nand2_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11054_ _164_\[22\] _01217_ _04627_ net50 _01423_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__o221a_1
X_10005_ _01292_ _04316_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__nor2_1
XFILLER_92_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11956_ _05946_ _05951_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__or2_1
XFILLER_44_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10907_ _164_\[4\] _167_\[4\] _05064_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__mux2_1
X_11887_ _01361_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__clkbuf_4
X_13626_ clknet_leaf_51_clk _00845_ VGND VGND VPWR VPWR _140_\[26\] sky130_fd_sc_hd__dfxtp_2
X_10838_ _04636_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__clkbuf_4
X_13557_ clknet_leaf_73_clk _00776_ VGND VGND VPWR VPWR _149_\[21\] sky130_fd_sc_hd__dfxtp_1
X_10769_ _04971_ _04978_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__or2_1
XFILLER_118_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13488_ clknet_leaf_50_clk _00707_ VGND VGND VPWR VPWR _158_\[6\] sky130_fd_sc_hd__dfxtp_1
X_12508_ _06290_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12439_ _06254_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07980_ _02513_ _02514_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__xnor2_1
X_06931_ _176_\[10\] _240_\[10\] _01449_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__mux2_1
XFILLER_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09650_ _04038_ _04039_ _04041_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__a21oi_1
X_06862_ _179_\[23\] _01301_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__or2_1
XFILLER_83_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08601_ _03023_ _03024_ _03030_ _01520_ _01439_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__o221a_1
X_09581_ _01278_ _03873_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__nor2_2
X_06793_ _246_\[5\] _01422_ _01425_ _01447_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__o211a_1
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08532_ _02947_ _02948_ _02963_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__o21a_1
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08463_ _02895_ _02876_ _02896_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__o21a_1
XFILLER_51_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07414_ _182_\[9\] _01632_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__nand2_1
XFILLER_51_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08394_ net49 _02798_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__or2_1
XFILLER_23_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07345_ _01868_ _01894_ _01900_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_30_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
X_07276_ _01806_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__inv_2
X_09015_ _03428_ _03431_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__nand2_1
XFILLER_105_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09917_ _142_\[16\] _04298_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_97_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_16
X_09848_ _04087_ _03958_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__or2_1
XFILLER_74_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _03910_ _04166_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__or2_1
XFILLER_100_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _140_\[18\] _05821_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__xnor2_1
X_12790_ _06438_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__clkbuf_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _152_\[2\] _05757_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__or2_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _116_\[25\] _05687_ _05677_ _116_\[24\] VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__o211a_1
XFILLER_53_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10623_ _176_\[15\] _04678_ _04627_ _173_\[15\] _02833_ VGND VGND VPWR VPWR _04878_
+ sky130_fd_sc_hd__o221a_1
XFILLER_41_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13411_ clknet_leaf_126_clk _00630_ VGND VGND VPWR VPWR _167_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
X_13342_ clknet_leaf_10_clk _00561_ VGND VGND VPWR VPWR _173_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10554_ _01213_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__clkbuf_4
XFILLER_139_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10485_ _04766_ _04781_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__or2_1
X_13273_ clknet_leaf_25_clk _00492_ VGND VGND VPWR VPWR _179_\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_142_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12224_ _06141_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12155_ _06105_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__clkbuf_1
X_11106_ _158_\[4\] _01254_ _05194_ _05196_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__o31a_1
XFILLER_111_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12086_ _06069_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_88_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_16
X_11037_ net42 _04848_ _05163_ _01436_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__a211o_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12988_ clknet_leaf_13_clk _00207_ VGND VGND VPWR VPWR _243_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11939_ net11 _05742_ _05938_ _05939_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__o22a_1
XFILLER_33_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13609_ clknet_leaf_52_clk _00828_ VGND VGND VPWR VPWR _140_\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_119_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07130_ _237_\[28\] VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_12_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07061_ _240_\[12\] _01601_ _01598_ _01644_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__o211a_1
XFILLER_145_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_79_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_16
X_07963_ _02497_ _02498_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__nor2_1
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09702_ _04047_ _04072_ _04092_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06914_ _176_\[5\] _01531_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__or2_1
XFILLER_68_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07894_ _02430_ _02431_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__xnor2_1
X_09633_ _03886_ _04025_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__nor2_1
XFILLER_110_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06845_ _243_\[18\] _01438_ _01486_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09564_ _01277_ _01282_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__nand2_2
XFILLER_55_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06776_ _01426_ _01433_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__nand2_1
X_08515_ _02919_ _02921_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__nor2_1
X_09495_ _03892_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__buf_2
X_08446_ _228_\[0\] _231_\[0\] _02768_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__a21o_1
XFILLER_24_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08377_ _228_\[17\] _02775_ _02810_ _02826_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__a211o_1
XFILLER_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07328_ _01623_ _01827_ _01693_ _01885_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__a211o_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07259_ _01802_ _01818_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__xor2_1
XFILLER_133_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10270_ _01305_ _01338_ _04624_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__or3_2
XFILLER_3_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13960_ clknet_leaf_71_clk _01179_ VGND VGND VPWR VPWR _118_\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12911_ clknet_leaf_74_clk _00135_ VGND VGND VPWR VPWR _116_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13891_ clknet_leaf_64_clk _01110_ VGND VGND VPWR VPWR _122_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12842_ _06465_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__clkbuf_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _06429_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__clkbuf_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _140_\[19\] _05743_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__xnor2_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _05665_ _05667_ _05672_ _05682_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__o31a_1
X_10606_ _173_\[9\] _04849_ _04866_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__a21bo_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11586_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__inv_2
X_13325_ clknet_leaf_22_clk _00544_ VGND VGND VPWR VPWR _173_\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_6_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10537_ _04671_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13256_ clknet_leaf_28_clk _00475_ VGND VGND VPWR VPWR _179_\[2\] sky130_fd_sc_hd__dfxtp_1
X_10468_ _176_\[1\] _179_\[1\] _04743_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__mux2_1
X_12207_ _06132_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13187_ clknet_leaf_33_clk _00406_ _00108_ VGND VGND VPWR VPWR _195_\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_111_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10399_ _04712_ _04719_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__or2_1
X_12138_ _06096_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12069_ _06058_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_1_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
X_06630_ _099_ _01295_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__nand2_1
XFILLER_92_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06561_ _01252_ _01269_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__or2_1
XFILLER_80_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06492_ _392_\[1\] _392_\[0\] VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__or2_2
X_09280_ _03651_ _03670_ _03688_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__o21ai_1
X_08300_ _231_\[31\] _02706_ _02765_ _02767_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__o211a_1
XFILLER_21_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08231_ _231_\[11\] _02706_ _02695_ _02718_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__o211a_1
XFILLER_118_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08162_ _167_\[24\] _02652_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__or2_1
XFILLER_118_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07113_ _173_\[24\] _01646_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__or2_1
X_08093_ _231_\[4\] _02611_ _01695_ _02619_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__o211a_1
XFILLER_134_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07044_ _240_\[8\] _01601_ _01598_ _01631_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__o211a_1
XFILLER_133_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08995_ _02835_ _02794_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07946_ _02473_ _02475_ _02472_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__o21a_1
XFILLER_28_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07877_ _02414_ _02415_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__or2_2
XFILLER_55_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09616_ _01280_ _03875_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__nor2b_4
X_06828_ _246_\[14\] _01407_ _01460_ _01473_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__a211o_1
XFILLER_83_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09547_ _03920_ _03942_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__or2_1
X_06759_ _01418_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__buf_4
X_09478_ _195_\[3\] _03875_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__nor2_4
XFILLER_51_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08429_ _02865_ _01801_ _02824_ _02866_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__o211a_1
XFILLER_11_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11440_ _05477_ _05481_ _05489_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11371_ _149_\[24\] _132_\[24\] _05429_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__a21o_1
X_10322_ _182_\[21\] _04654_ _04642_ _04650_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__a31o_1
X_13110_ clknet_leaf_118_clk _00329_ VGND VGND VPWR VPWR _231_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13041_ clknet_leaf_110_clk _00260_ VGND VGND VPWR VPWR _237_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10253_ _04613_ _04619_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10184_ _04529_ _04550_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__nand2_1
XFILLER_79_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13943_ clknet_leaf_91_clk _01162_ VGND VGND VPWR VPWR _120_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13874_ clknet_leaf_96_clk _01093_ VGND VGND VPWR VPWR _124_\[18\] sky130_fd_sc_hd__dfxtp_1
X_12825_ _06456_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12756_ _06420_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _06384_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__clkbuf_1
X_11707_ _149_\[29\] _05729_ _05625_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__mux2_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11638_ _05665_ _05667_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__xor2_1
X_11569_ _05604_ _05605_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__xnor2_1
X_13308_ clknet_leaf_4_clk _00527_ VGND VGND VPWR VPWR _176_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13239_ clknet_leaf_25_clk _00458_ VGND VGND VPWR VPWR _182_\[17\] sky130_fd_sc_hd__dfxtp_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08780_ _03201_ _03203_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__xnor2_1
X_07800_ _02339_ _02340_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__and2_1
XFILLER_85_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07731_ _02248_ _02250_ _02273_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__o21ba_1
XFILLER_77_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07662_ _01684_ _01638_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__xnor2_2
X_06613_ _01315_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__clkbuf_4
X_07593_ _01444_ _02140_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__nand2_1
X_09401_ _170_\[29\] _02865_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__nand2_1
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06544_ _01249_ _01252_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__nor2_2
XFILLER_111_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09332_ _03689_ _03728_ _03738_ _03694_ _03729_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__o221a_1
XFILLER_33_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09263_ _185_\[25\] _03644_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nand2_1
XFILLER_21_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09194_ _170_\[23\] _02846_ _03604_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__a21oi_1
X_08214_ _01799_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__buf_2
X_08145_ _167_\[19\] _02652_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__or2_1
XFILLER_112_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08076_ _01355_ _02603_ _02607_ _02355_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__a211o_1
XFILLER_134_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07027_ _01615_ _01618_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__or2_1
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08978_ _03380_ _03381_ _03394_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__nor3_1
XFILLER_29_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07929_ _02396_ _02436_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__nand2_1
XFILLER_90_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10940_ net40 _05068_ _05100_ _05086_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__a211o_1
XFILLER_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12610_ _128_\[30\] _126_\[30\] _06335_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__mux2_1
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10871_ _05028_ _05051_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__or2_1
X_13590_ clknet_leaf_48_clk _00809_ VGND VGND VPWR VPWR _142_\[22\] sky130_fd_sc_hd__dfxtp_2
XFILLER_129_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12541_ _130_\[29\] _128_\[29\] _06302_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__mux2_1
XFILLER_61_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12472_ _132_\[28\] _130_\[28\] _06269_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__mux2_1
XFILLER_61_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11423_ _118_\[7\] _118_\[3\] VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 _03667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11354_ _152_\[22\] _05262_ _05413_ _05415_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__a22o_1
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10305_ _182_\[13\] _04634_ _04657_ _04649_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__o211a_1
X_11285_ _149_\[14\] _132_\[14\] VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__nand2_1
X_10236_ _04582_ _04585_ _04603_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__o21ba_1
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13024_ clknet_leaf_17_clk _00243_ VGND VGND VPWR VPWR _237_\[0\] sky130_fd_sc_hd__dfxtp_4
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10167_ _246_\[27\] _01316_ _04409_ _243_\[27\] _01507_ VGND VGND VPWR VPWR _04538_
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10098_ _142_\[24\] _04471_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__and2_1
XFILLER_94_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13926_ clknet_leaf_70_clk _01145_ VGND VGND VPWR VPWR _120_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13857_ clknet_leaf_69_clk _01076_ VGND VGND VPWR VPWR _124_\[1\] sky130_fd_sc_hd__dfxtp_1
X_13788_ clknet_leaf_68_clk _01007_ VGND VGND VPWR VPWR _130_\[28\] sky130_fd_sc_hd__dfxtp_1
X_12808_ _06447_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12739_ _06411_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__clkbuf_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09950_ _04308_ _04311_ _04329_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__a21boi_1
XFILLER_89_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08901_ _03281_ _03283_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__nor2_1
X_09881_ _142_\[13\] _04228_ _04240_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08832_ _02855_ _03253_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__xnor2_2
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _03170_ _03171_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__nand2_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07714_ _02218_ _02238_ _02256_ _01269_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__a31o_1
XFILLER_38_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08694_ _03119_ _03120_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__nor2_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07645_ _02189_ _02190_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__or2_1
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07576_ _02089_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__inv_2
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06527_ _01235_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__buf_2
XFILLER_80_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09315_ _03679_ _03708_ _03721_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__and3_1
X_09246_ _03653_ _03655_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09177_ _03587_ _03588_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__and2b_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08128_ _231_\[14\] _02611_ _02641_ _02644_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__o211a_1
X_08059_ _01704_ _02564_ _02178_ _02591_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__a211o_1
XFILLER_122_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput46 net46 VGND VGND VPWR VPWR dout[19] sky130_fd_sc_hd__buf_2
X_11070_ _04638_ _05183_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__or2_1
Xoutput57 net57 VGND VGND VPWR VPWR dout[29] sky130_fd_sc_hd__buf_2
X_10021_ _04345_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__inv_2
Xoutput68 net68 VGND VGND VPWR VPWR dst_write sky130_fd_sc_hd__buf_2
XFILLER_103_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11972_ _05955_ _05961_ _05969_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__o21bai_1
X_13711_ clknet_leaf_78_clk _00930_ VGND VGND VPWR VPWR _134_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10923_ net66 _05048_ _05088_ _05067_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__o211a_1
XFILLER_17_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13642_ clknet_leaf_48_clk _00861_ VGND VGND VPWR VPWR _138_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10854_ _05028_ _05039_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__or2_1
XFILLER_32_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13573_ clknet_leaf_53_clk _00792_ VGND VGND VPWR VPWR _142_\[5\] sky130_fd_sc_hd__dfxtp_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ _130_\[21\] _128_\[21\] _06291_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__mux2_1
X_10785_ _164_\[0\] _04983_ _04990_ _04939_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__o211a_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12455_ _132_\[20\] _130_\[20\] _06258_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__mux2_1
X_11406_ _05458_ _05459_ _05460_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__and3_1
X_12386_ _132_\[19\] _134_\[19\] _06219_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__mux2_1
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11337_ _152_\[20\] _01368_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__and2_1
XFILLER_141_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11268_ _05340_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__clkbuf_1
X_11199_ _149_\[3\] _132_\[3\] VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__nor2_1
X_10219_ _04558_ _04573_ _04587_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__o21ba_1
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13007_ clknet_leaf_18_clk _00226_ VGND VGND VPWR VPWR _240_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13909_ clknet_leaf_93_clk _01128_ VGND VGND VPWR VPWR _122_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07430_ _01954_ _01975_ _01981_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__nand3_1
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07361_ _182_\[8\] _01629_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__nand2_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09100_ _03486_ _03488_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__or2b_1
X_07292_ _01802_ _01818_ _01816_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__a21oi_1
X_09031_ _185_\[18\] _03413_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__nand2_1
XFILLER_117_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09933_ _01243_ _01281_ _03960_ _03888_ _04132_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__a32o_1
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09864_ _185_\[13\] _04150_ _04175_ _04248_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__o211a_1
XFILLER_100_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08815_ _03173_ _03237_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__or2_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _03933_ _04181_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__nor2_1
XFILLER_85_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08746_ _03147_ _03148_ _03149_ _03146_ _03144_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__o32ai_2
XFILLER_54_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _185_\[8\] _03103_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__xnor2_2
XFILLER_54_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07628_ _02173_ _02174_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__nor2_2
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07559_ _02106_ _02107_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__nand2_1
X_10570_ _176_\[30\] _179_\[30\] _04830_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__mux2_1
XFILLER_127_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09229_ _03622_ _03624_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__and2b_1
XFILLER_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12240_ _138_\[14\] _136_\[14\] _06145_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__mux2_1
XFILLER_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12171_ _140_\[13\] _138_\[13\] _06112_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__mux2_1
XFILLER_5_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11122_ _158_\[7\] _01256_ _158_\[8\] VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11053_ net49 _04628_ _05173_ _05117_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__o211a_1
X_10004_ _04076_ _04104_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__nand2_1
XFILLER_67_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11955_ _05954_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10906_ net61 _05048_ _05076_ _05067_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__o211a_1
X_13625_ clknet_leaf_49_clk _00844_ VGND VGND VPWR VPWR _140_\[25\] sky130_fd_sc_hd__dfxtp_2
X_11886_ net6 _05891_ _05852_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__mux2_1
X_10837_ _164_\[15\] _05025_ _05027_ _05001_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__a211o_1
X_13556_ clknet_leaf_73_clk _00775_ VGND VGND VPWR VPWR _149_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10768_ _170_\[28\] _173_\[28\] _04936_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__mux2_1
XFILLER_13_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13487_ clknet_leaf_36_clk _00706_ VGND VGND VPWR VPWR _158_\[5\] sky130_fd_sc_hd__dfxtp_1
X_12507_ _130_\[13\] _128_\[13\] _06280_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__mux2_1
X_12438_ _132_\[12\] _130_\[12\] _06247_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__mux2_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10699_ _167_\[7\] _04925_ _04929_ _04891_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__o211a_1
XFILLER_141_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12369_ _132_\[11\] _134_\[11\] _06208_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__mux2_1
XFILLER_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06930_ _01421_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__buf_2
X_06861_ _246_\[22\] _01496_ _01460_ _01498_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__a211o_1
XFILLER_94_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08600_ _03029_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__inv_2
X_09580_ _142_\[3\] _03974_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__xnor2_1
X_06792_ _01444_ _01446_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__nand2_1
XFILLER_83_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08531_ _02960_ _02962_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08462_ _185_\[0\] _02875_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__nand2_1
X_07413_ _182_\[9\] _01632_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__or2_1
XFILLER_50_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08393_ _225_\[21\] VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__buf_4
X_07344_ _01868_ _01894_ _01900_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07275_ _01813_ _01814_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__and2b_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09014_ _03368_ _03429_ _03430_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__o21bai_1
XFILLER_117_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09916_ _246_\[16\] _01315_ _04129_ _243_\[16\] _01477_ VGND VGND VPWR VPWR _04298_
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09847_ _01281_ _04231_ _03908_ _01231_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__a211oi_1
XFILLER_100_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _04163_ _04164_ _04165_ _03872_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__o22a_1
XFILLER_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _01408_ _03153_ _03154_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__or3_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _152_\[2\] _05757_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__nand2_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _05680_ _05688_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__or2_1
X_10622_ _04853_ _04876_ _04877_ _04839_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__a211o_1
XFILLER_41_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13410_ clknet_leaf_126_clk _00629_ VGND VGND VPWR VPWR _167_\[28\] sky130_fd_sc_hd__dfxtp_2
X_10553_ _173_\[25\] _04774_ _04829_ _04777_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__a211o_1
X_13341_ clknet_leaf_4_clk _00560_ VGND VGND VPWR VPWR _173_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10484_ _176_\[5\] _179_\[5\] _04743_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__mux2_1
X_13272_ clknet_leaf_25_clk _00491_ VGND VGND VPWR VPWR _179_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12223_ _138_\[6\] _136_\[6\] _06134_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__mux2_1
XFILLER_142_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12154_ _140_\[5\] _138_\[5\] _06101_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__mux2_1
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11105_ net5 _05196_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__nor2_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12085_ _140_\[4\] _142_\[4\] _06068_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__mux2_1
XFILLER_96_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11036_ _164_\[15\] _04872_ _04633_ _05162_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__o211a_1
XFILLER_92_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12987_ clknet_leaf_13_clk _00206_ VGND VGND VPWR VPWR _243_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11938_ _05936_ _05937_ _05785_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__o21ai_1
XFILLER_72_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11869_ _152_\[13\] _05875_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__nand2_1
X_13608_ clknet_leaf_53_clk _00827_ VGND VGND VPWR VPWR _140_\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13539_ clknet_leaf_65_clk _00758_ VGND VGND VPWR VPWR _149_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07060_ _01615_ _01643_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__or2_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09701_ _04074_ _04091_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__xor2_1
X_07962_ _02457_ _02484_ _02496_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__o21a_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06913_ _01495_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07893_ _243_\[25\] _240_\[25\] _01687_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__mux2_4
X_09632_ _03903_ _03880_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__nand2_1
X_06844_ _179_\[18\] _01300_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__or2_1
XFILLER_95_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09563_ _03957_ _03958_ _195_\[4\] VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__a21oi_1
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06775_ _243_\[2\] _01428_ _01432_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__o21ai_1
X_08514_ _02945_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__inv_2
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09494_ _01240_ _03890_ _03891_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__and3_1
XFILLER_70_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08445_ _02878_ _02879_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__nand2_1
X_08376_ _02823_ _02791_ _02824_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__o211a_1
XFILLER_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07327_ _01856_ _01863_ _01883_ _01884_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__a211oi_1
XFILLER_139_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07258_ _01816_ _01817_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__nor2_1
XFILLER_136_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07189_ _01746_ _01750_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13890_ clknet_leaf_64_clk _01109_ VGND VGND VPWR VPWR _122_\[2\] sky130_fd_sc_hd__dfxtp_1
X_12910_ clknet_leaf_89_clk _00134_ VGND VGND VPWR VPWR _116_\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12841_ _118_\[12\] _120_\[12\] _06462_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__mux2_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12772_ _122_\[11\] _120_\[11\] _06423_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__mux2_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _140_\[17\] _140_\[10\] VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__xnor2_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _116_\[23\] _05671_ _05681_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__o21ai_1
XFILLER_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10605_ _04864_ _04678_ _01971_ _04865_ _02833_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__o221a_1
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11585_ _116_\[17\] _05618_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__nor2_1
X_13324_ clknet_leaf_22_clk _00543_ VGND VGND VPWR VPWR _173_\[6\] sky130_fd_sc_hd__dfxtp_2
X_10536_ _173_\[20\] _04780_ _04817_ _04785_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__o211a_1
XFILLER_6_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10467_ _173_\[0\] _04735_ _04768_ _04740_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__o211a_1
X_13255_ clknet_leaf_24_clk _00474_ VGND VGND VPWR VPWR _179_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12206_ _140_\[30\] _138_\[30\] _06123_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__mux2_1
XFILLER_108_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13186_ clknet_leaf_33_clk _00405_ _00107_ VGND VGND VPWR VPWR _195_\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_96_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10398_ _179_\[13\] _182_\[13\] _04693_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__mux2_1
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12137_ _140_\[29\] _142_\[29\] _06090_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__mux2_1
XFILLER_111_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12068_ _142_\[30\] _06057_ _06005_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__mux2_1
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11019_ _164_\[9\] net68 _03133_ _04692_ _01417_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__a221o_1
XFILLER_92_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06560_ _01268_ _01251_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__nor2_8
XFILLER_52_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08230_ _02686_ _02717_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__or2_1
XFILLER_60_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08161_ _234_\[23\] _02659_ _02636_ _02668_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__o211a_1
XFILLER_118_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07112_ _237_\[24\] VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__buf_4
X_08092_ _167_\[4\] _02616_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__or2_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07043_ _01615_ _01630_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__or2_1
XFILLER_142_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08994_ _03391_ _03393_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__and2b_1
X_07945_ _02479_ _02480_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__or2b_1
XFILLER_29_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09615_ _04002_ _03957_ _03903_ _03899_ _01235_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__a311o_1
XFILLER_141_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07876_ _02405_ _02406_ _02413_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06827_ _243_\[14\] _01438_ _01461_ _01472_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__o211a_1
XFILLER_83_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09546_ _03920_ _03942_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__nand2_1
X_06758_ _01417_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__clkbuf_4
XFILLER_36_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09477_ _03874_ _01282_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__nor2_4
XFILLER_24_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06689_ _01376_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08428_ net57 _01519_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__or2_1
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08359_ _02811_ _02791_ _02760_ _02812_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__o211a_1
XFILLER_109_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11370_ _05421_ _05423_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__and2b_1
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10321_ _182_\[20\] _04663_ _04666_ _04649_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__o211a_1
XFILLER_3_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13040_ clknet_leaf_83_clk _00259_ VGND VGND VPWR VPWR _237_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10252_ _142_\[31\] _04618_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10183_ _185_\[27\] _03870_ _03864_ _04553_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__o211a_1
XFILLER_78_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13942_ clknet_leaf_96_clk _01161_ VGND VGND VPWR VPWR _120_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13873_ clknet_leaf_95_clk _01092_ VGND VGND VPWR VPWR _124_\[17\] sky130_fd_sc_hd__dfxtp_1
X_12824_ _118_\[4\] _120_\[4\] _06451_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__mux2_1
XFILLER_74_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12755_ _122_\[3\] _120_\[3\] _06412_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__mux2_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11706_ _05727_ _05728_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__xnor2_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12686_ _124_\[2\] _122_\[2\] _06379_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__mux2_1
XFILLER_91_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11637_ _05639_ _05648_ _05649_ _05658_ _05666_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__o41a_1
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11568_ _05595_ _05597_ _05593_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__o21ai_1
XFILLER_7_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10519_ _173_\[15\] _04780_ _04805_ _04785_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__o211a_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13307_ clknet_leaf_4_clk _00526_ VGND VGND VPWR VPWR _176_\[21\] sky130_fd_sc_hd__dfxtp_1
X_11499_ _116_\[8\] _05541_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__or2_1
X_13238_ clknet_leaf_25_clk _00457_ VGND VGND VPWR VPWR _182_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13169_ clknet_leaf_105_clk _00388_ VGND VGND VPWR VPWR _225_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07730_ _02251_ _02252_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__and2b_1
XFILLER_38_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07661_ _02205_ _02187_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__or2_1
XFILLER_37_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06612_ _01314_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__buf_2
XFILLER_80_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07592_ _02134_ _02139_ _01427_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__mux2_1
XFILLER_53_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09400_ _170_\[29\] _02865_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__or2_1
X_06543_ _01250_ _01251_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__nor2_2
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09331_ _03691_ _03730_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__nand2_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09262_ _02431_ _03649_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__nand2_1
XFILLER_21_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08213_ _231_\[6\] _02690_ _02664_ _02705_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__a211o_1
X_09193_ _170_\[23\] _02846_ _02842_ _170_\[22\] _03603_ VGND VGND VPWR VPWR _03604_
+ sky130_fd_sc_hd__o221a_1
X_08144_ _234_\[18\] _02646_ _02629_ _02656_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__a211o_1
XFILLER_119_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08075_ _01778_ _02606_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__nor2_1
X_07026_ _173_\[4\] _01616_ _01617_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__mux2_1
XFILLER_103_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08977_ _03380_ _03381_ _03394_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07928_ _02463_ _02464_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__and2_1
X_07859_ _02339_ _02373_ _02397_ _02344_ _02374_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__o221a_1
XFILLER_28_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10870_ _167_\[25\] _170_\[25\] _04995_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__mux2_1
X_09529_ _03883_ _03925_ _01240_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__mux2_1
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12540_ _06307_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12471_ _06271_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11422_ _05474_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11353_ _05352_ _05414_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__nor2_1
XFILLER_106_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10304_ _179_\[13\] _04646_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__or2_1
X_11284_ _149_\[14\] _132_\[14\] VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__or2_1
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10235_ _04600_ _04602_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__xnor2_1
X_13023_ clknet_leaf_13_clk _00242_ VGND VGND VPWR VPWR _240_\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10166_ _04529_ _04534_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__nand2_1
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10097_ _246_\[24\] _01315_ _04409_ _243_\[24\] _01501_ VGND VGND VPWR VPWR _04471_
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13925_ clknet_leaf_70_clk _01144_ VGND VGND VPWR VPWR _120_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13856_ clknet_leaf_64_clk _01075_ VGND VGND VPWR VPWR _124_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12807_ _122_\[28\] _120_\[28\] _01367_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__mux2_1
X_13787_ clknet_leaf_68_clk _01006_ VGND VGND VPWR VPWR _130_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10999_ net36 _164_\[0\] _01215_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__mux2_1
X_12738_ _124_\[27\] _122_\[27\] _06401_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__mux2_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ _126_\[26\] _124_\[26\] _06368_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__mux2_1
XFILLER_129_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09880_ _04262_ _04263_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__or2_1
XFILLER_98_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08900_ _02127_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__xnor2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08831_ _02817_ _225_\[3\] VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__xnor2_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _02801_ _03032_ _02861_ _03186_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__a211o_1
X_07713_ _02218_ _02238_ _02256_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__a21oi_1
X_08693_ _170_\[8\] _02794_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__and2_1
XFILLER_38_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07644_ _02153_ _02155_ _02188_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__and3_1
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07575_ _02121_ _02122_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__nand2_1
XFILLER_53_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06526_ _01234_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__buf_2
X_09314_ _03679_ _03708_ _03721_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__a21oi_1
X_09245_ _228_\[25\] _231_\[25\] _03654_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__o21a_1
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09176_ _03571_ _03572_ _03586_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__o21ai_1
XFILLER_119_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08127_ _167_\[14\] _02616_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__or2_1
XFILLER_135_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08058_ _01520_ _02570_ _02590_ _02202_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__o211a_1
Xoutput47 net47 VGND VGND VPWR VPWR dout[1] sky130_fd_sc_hd__buf_2
XFILLER_122_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07009_ _237_\[1\] VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__clkbuf_4
Xoutput36 net36 VGND VGND VPWR VPWR dout[0] sky130_fd_sc_hd__buf_2
Xoutput58 net58 VGND VGND VPWR VPWR dout[2] sky130_fd_sc_hd__buf_2
Xoutput69 net69 VGND VGND VPWR VPWR src_read sky130_fd_sc_hd__buf_2
X_10020_ _04295_ _04296_ _04397_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__a21o_1
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11971_ _05944_ _05960_ _05959_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13710_ clknet_leaf_78_clk _00929_ VGND VGND VPWR VPWR _134_\[14\] sky130_fd_sc_hd__dfxtp_1
X_10922_ _05079_ _05087_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__or2_1
XFILLER_29_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13641_ clknet_leaf_54_clk _00860_ VGND VGND VPWR VPWR _138_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_776 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10853_ _167_\[20\] _170_\[20\] _04995_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__mux2_1
XFILLER_32_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13572_ clknet_leaf_52_clk _00791_ VGND VGND VPWR VPWR _142_\[4\] sky130_fd_sc_hd__dfxtp_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10784_ _04971_ _04989_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__or2_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _06298_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__clkbuf_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12454_ _06262_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11405_ _05452_ _05454_ _05453_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__a21boi_1
X_12385_ _06226_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11336_ _05381_ _05386_ _05389_ _05397_ _05388_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__a311o_2
XFILLER_113_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11267_ _152_\[11\] _05339_ _05318_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__mux2_1
X_13006_ clknet_leaf_14_clk _00225_ VGND VGND VPWR VPWR _240_\[14\] sky130_fd_sc_hd__dfxtp_1
X_10218_ _04585_ _04586_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__or2_1
X_11198_ _05263_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__buf_4
X_10149_ _01281_ _03876_ _04520_ _04210_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__a211o_1
XFILLER_121_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13908_ clknet_leaf_92_clk _01127_ VGND VGND VPWR VPWR _122_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13839_ clknet_leaf_95_clk _01058_ VGND VGND VPWR VPWR _126_\[15\] sky130_fd_sc_hd__dfxtp_1
X_07360_ _182_\[8\] _01629_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__or2_1
XFILLER_62_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07291_ _01811_ _01834_ _01848_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__o21a_1
X_09030_ _02242_ _03445_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09932_ _185_\[16\] _04150_ _04175_ _04313_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__o211a_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09863_ _03945_ _04246_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__or3_1
XFILLER_112_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _03898_ _03893_ _03876_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__a21oi_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08814_ _03205_ _03206_ _03172_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__nand3b_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _03167_ _03169_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08676_ _02868_ _03102_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__xnor2_4
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07627_ _02170_ _02172_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__and2_1
X_07558_ _182_\[14\] _01650_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__nand2_1
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06509_ _01218_ _01219_ _01221_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__o21a_1
XFILLER_42_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07489_ _01681_ _02039_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09228_ _03620_ _03621_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__and2b_1
XFILLER_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09159_ _03555_ _03557_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__and2b_1
XFILLER_107_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12170_ _06113_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11121_ _158_\[7\] _05193_ _05218_ _05191_ _05219_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__a221o_1
XFILLER_122_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11052_ _04638_ _05172_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__or2_1
X_10003_ _04379_ _04380_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__or2_1
XFILLER_77_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11954_ _142_\[20\] _05953_ _05893_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__mux2_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11885_ _05888_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__xor2_1
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10905_ _05028_ _05075_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__or2_1
X_13624_ clknet_leaf_50_clk _00843_ VGND VGND VPWR VPWR _140_\[24\] sky130_fd_sc_hd__dfxtp_2
XFILLER_72_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10836_ _167_\[15\] _05022_ _05009_ _05026_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__o211a_1
XFILLER_32_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13555_ clknet_leaf_74_clk _00774_ VGND VGND VPWR VPWR _149_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10767_ _167_\[27\] _04925_ _04977_ _04939_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__o211a_1
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13486_ clknet_leaf_36_clk _00705_ VGND VGND VPWR VPWR _158_\[4\] sky130_fd_sc_hd__dfxtp_1
X_12506_ _06289_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10698_ _04888_ _04928_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__or2_1
XFILLER_145_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12437_ _06253_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12368_ _06217_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12299_ _136_\[10\] _134_\[10\] _06178_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__mux2_1
X_11319_ _05383_ _05384_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__nand2_1
XFILLER_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06860_ _243_\[22\] _01474_ _01461_ _01497_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__o211a_1
XFILLER_68_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06791_ _243_\[5\] _01428_ _01445_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__o21ai_1
XFILLER_82_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08530_ _228_\[3\] _231_\[3\] _02961_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__o21a_1
X_08461_ _01714_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__inv_2
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07412_ _01949_ _01964_ _01354_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__o21a_1
X_08392_ _01406_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07343_ _01896_ _01899_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__xor2_1
XFILLER_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07274_ _01832_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__inv_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09013_ _03400_ _03395_ _03396_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__a21oi_1
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09915_ _04277_ _04285_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__nor2_1
X_09846_ _01242_ _04230_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__or2_1
XFILLER_113_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _03884_ _03898_ _03873_ _04006_ _04051_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__a32o_1
XFILLER_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06989_ _176_\[27\] _01580_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__or2_1
XFILLER_39_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08728_ _03134_ _03135_ _03152_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _03048_ _03049_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__nand2_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _05694_ _05695_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__nand2_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10621_ _02111_ _04631_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__nor2_1
XFILLER_139_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10552_ _176_\[25\] _04771_ _04806_ _04828_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__o211a_1
X_13340_ clknet_leaf_4_clk _00559_ VGND VGND VPWR VPWR _173_\[22\] sky130_fd_sc_hd__dfxtp_1
X_13271_ clknet_leaf_7_clk _00490_ VGND VGND VPWR VPWR _179_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12222_ _06140_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__clkbuf_1
X_10483_ _04671_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12153_ _06104_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12084_ _06004_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__clkbuf_4
X_11104_ net4 _05202_ _05193_ _158_\[3\] _05206_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__a221o_1
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11035_ _03338_ _04681_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__nand2_1
XFILLER_77_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12986_ clknet_leaf_13_clk _00205_ VGND VGND VPWR VPWR _243_\[26\] sky130_fd_sc_hd__dfxtp_1
X_11937_ _05936_ _05937_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__and2_1
X_11868_ _140_\[23\] _05874_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__xnor2_1
X_13607_ clknet_leaf_53_clk _00826_ VGND VGND VPWR VPWR _140_\[7\] sky130_fd_sc_hd__dfxtp_1
X_11799_ _140_\[24\] _140_\[26\] VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10819_ _04971_ _05014_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__or2_1
X_13538_ clknet_leaf_66_clk _00757_ VGND VGND VPWR VPWR _149_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13469_ clknet_leaf_129_clk _00688_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfxtp_1
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07961_ _02457_ _02484_ _02496_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__nor3_1
X_09700_ _01231_ _04079_ _04084_ _04090_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__a31o_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06912_ _243_\[4\] _01485_ _01481_ _01535_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__o211a_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07892_ _02428_ _02429_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__or2_1
X_09631_ _142_\[5\] _04023_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06843_ _01421_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__clkbuf_4
XFILLER_95_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09562_ _01277_ _195_\[3\] VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__and2b_1
X_06774_ _179_\[2\] _01268_ _01251_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__or3_1
XFILLER_83_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08513_ _02942_ _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__xor2_1
X_09493_ _03874_ _195_\[0\] VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__or2b_1
XFILLER_91_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08444_ _01719_ _02877_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__or2_1
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08375_ net44 _02798_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__or2_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07326_ _01405_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__clkbuf_8
XFILLER_32_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07257_ _01786_ _01803_ _01815_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__nor3_1
XFILLER_145_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07188_ _01748_ _01749_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__nor2_1
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09829_ _04002_ _04005_ _03933_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__a21o_1
XFILLER_86_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12840_ _06464_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__clkbuf_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12771_ _06428_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__clkbuf_1
X_11722_ _01358_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__buf_4
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _116_\[22\] _05662_ _05671_ _116_\[23\] VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__a22o_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10604_ _04625_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__buf_4
XFILLER_127_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13323_ clknet_leaf_23_clk _00542_ VGND VGND VPWR VPWR _173_\[5\] sky130_fd_sc_hd__dfxtp_1
X_11584_ _116_\[17\] _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__nand2_1
X_10535_ _04809_ _04816_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__or2_1
XFILLER_142_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13254_ clknet_leaf_24_clk _00473_ VGND VGND VPWR VPWR _179_\[0\] sky130_fd_sc_hd__dfxtp_1
X_10466_ _04766_ _04767_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__or2_1
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13185_ clknet_leaf_33_clk _00404_ _00106_ VGND VGND VPWR VPWR _195_\[1\] sky130_fd_sc_hd__dfrtp_2
X_12205_ _06131_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12136_ _06095_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10397_ _176_\[12\] _04683_ _04718_ _01419_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__a211o_1
XFILLER_96_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12067_ _05742_ _06054_ _06055_ _06056_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__a31o_1
XFILLER_96_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11018_ _164_\[8\] _01218_ _03864_ _05151_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__o211a_1
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12969_ clknet_leaf_20_clk _00188_ VGND VGND VPWR VPWR _243_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08160_ _02625_ _02667_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__or2_1
X_07111_ _240_\[23\] _01660_ _01653_ _01683_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__o211a_1
X_08091_ _234_\[3\] _02564_ _02178_ _02618_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__a211o_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07042_ _173_\[8\] _01629_ _01617_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__mux2_1
XFILLER_133_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08993_ _03389_ _03390_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__nor2_1
X_07944_ _182_\[27\] _01694_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__nand2_1
XFILLER_68_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07875_ _02405_ _02406_ _02413_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__and3_1
XFILLER_56_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09614_ _03933_ _04001_ _04003_ _04007_ _01230_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__o221a_1
XFILLER_141_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06826_ _179_\[14\] _01300_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__or2_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09545_ _03922_ _03941_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06757_ _01416_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__buf_4
XFILLER_55_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_129_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_129_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_24_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09476_ _195_\[2\] VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__buf_2
X_06688_ _118_\[9\] _116_\[9\] _01370_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__mux2_1
X_08427_ _225_\[29\] VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__buf_4
XFILLER_24_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08358_ net40 _02798_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__or2_1
XFILLER_109_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07309_ _01707_ _01866_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__xnor2_2
X_08289_ _231_\[28\] _02730_ _02753_ _02759_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__a211o_1
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10320_ _179_\[20\] _04646_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__or2_1
X_10251_ _04210_ _04614_ _04615_ _04617_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__a31o_1
XFILLER_133_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10182_ _03945_ _04551_ _04552_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__or3_1
XFILLER_105_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13941_ clknet_leaf_93_clk _01160_ VGND VGND VPWR VPWR _120_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13872_ clknet_leaf_96_clk _01091_ VGND VGND VPWR VPWR _124_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12823_ _06455_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12754_ _06419_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__clkbuf_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11705_ _05715_ _05719_ _05713_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__o21ai_1
XFILLER_70_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12685_ _06383_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__clkbuf_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ _05646_ _05655_ _05656_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__a21o_1
X_11567_ _05602_ _05603_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__or2b_1
X_10518_ _04766_ _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__or2_1
XFILLER_7_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13306_ clknet_leaf_4_clk _00525_ VGND VGND VPWR VPWR _176_\[20\] sky130_fd_sc_hd__dfxtp_1
X_13237_ clknet_leaf_25_clk _00456_ VGND VGND VPWR VPWR _182_\[15\] sky130_fd_sc_hd__dfxtp_1
X_11498_ _116_\[8\] _05541_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__nand2_1
XFILLER_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10449_ _182_\[27\] _04746_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__or2_1
XFILLER_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13168_ clknet_leaf_105_clk _00387_ VGND VGND VPWR VPWR _225_\[16\] sky130_fd_sc_hd__dfxtp_1
X_12119_ _06086_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__clkbuf_1
X_13099_ clknet_leaf_106_clk _00318_ VGND VGND VPWR VPWR _231_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07660_ _02184_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__inv_2
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06611_ _01313_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__buf_2
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07591_ _02137_ _02138_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__xnor2_2
XFILLER_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06542_ _01207_ _01208_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__nand2_4
XFILLER_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09330_ _02858_ _03032_ _03309_ _03737_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__a211o_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09261_ _03653_ _03655_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__and2b_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08212_ _228_\[6\] _02698_ _02679_ _02704_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__o211a_1
X_09192_ _03509_ _03602_ _03540_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__a21o_1
XFILLER_21_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08143_ _231_\[18\] _02649_ _02641_ _02655_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__o211a_1
XFILLER_107_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08074_ _02604_ _02605_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__xnor2_2
X_07025_ _01518_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__clkbuf_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08976_ _03391_ _03393_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07927_ _02428_ _02449_ _02461_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__or3_1
XFILLER_29_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07858_ _02341_ _02375_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__nand2_1
X_06809_ _246_\[9\] _01422_ _01425_ _01459_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__o211a_1
XFILLER_44_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07789_ _02328_ _02329_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__nand2_1
X_09528_ _03924_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__buf_2
XFILLER_71_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09459_ _01856_ _03862_ _01884_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__a21oi_1
XFILLER_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12470_ _132_\[27\] _130_\[27\] _06269_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__mux2_1
XFILLER_8_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11421_ _152_\[31\] _05473_ _05439_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__mux2_1
X_11352_ _05395_ _05400_ _05403_ _05411_ _05402_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__a311oi_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10303_ _182_\[12\] _04634_ _04656_ _04649_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__o211a_1
X_11283_ _05351_ _05353_ _152_\[13\] _05262_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_140_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10234_ _142_\[30\] _04601_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__xor2_1
XFILLER_106_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13022_ clknet_leaf_11_clk _00241_ VGND VGND VPWR VPWR _240_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10165_ _03946_ _04535_ _04536_ _00105_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__o211a_1
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10096_ _185_\[23\] _03870_ _03864_ _04470_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__o211a_1
XFILLER_94_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13924_ clknet_leaf_70_clk _01143_ VGND VGND VPWR VPWR _120_\[4\] sky130_fd_sc_hd__dfxtp_1
X_13855_ clknet_leaf_65_clk _01074_ VGND VGND VPWR VPWR _126_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12806_ _06446_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13786_ clknet_leaf_68_clk _01005_ VGND VGND VPWR VPWR _130_\[26\] sky130_fd_sc_hd__dfxtp_1
X_10998_ net60 _05110_ _05140_ _05122_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__a211o_1
X_12737_ _06410_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__clkbuf_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _06374_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__clkbuf_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11619_ _05639_ _05649_ _05648_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12599_ _06338_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _03229_ _03232_ _03228_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__a21o_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08761_ _02380_ _03178_ _03185_ _02202_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__o211a_1
XFILLER_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07712_ _02254_ _02255_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__nor2_1
X_08692_ _170_\[8\] _02794_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__nor2_1
XFILLER_38_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07643_ _02153_ _02155_ _02188_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07574_ _02117_ _02120_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__nand2_1
X_09313_ _02495_ _03720_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06525_ _195_\[4\] VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__buf_2
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_16
X_09244_ _228_\[25\] _231_\[25\] _02852_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__a21o_1
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09175_ _03571_ _03572_ _03586_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__nor3_1
XFILLER_21_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08126_ _234_\[13\] _02564_ _02629_ _02643_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__a211o_1
X_08057_ _01408_ _02589_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__or2_1
Xoutput37 net37 VGND VGND VPWR VPWR dout[10] sky130_fd_sc_hd__buf_2
X_07008_ _240_\[0\] _01601_ _01598_ _01603_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__o211a_1
Xoutput48 net48 VGND VGND VPWR VPWR dout[20] sky130_fd_sc_hd__buf_2
Xoutput59 net59 VGND VGND VPWR VPWR dout[30] sky130_fd_sc_hd__buf_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08959_ _02380_ _03369_ _03377_ _01439_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__o211a_1
X_11970_ _05966_ _05967_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__nand2_1
XFILLER_57_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10921_ _164_\[8\] _167_\[8\] _05064_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__mux2_1
X_13640_ clknet_leaf_54_clk _00859_ VGND VGND VPWR VPWR _138_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10852_ _164_\[19\] _05025_ _05038_ _05035_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__a211o_1
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13571_ clknet_leaf_34_clk _00790_ VGND VGND VPWR VPWR _142_\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10783_ _167_\[0\] _170_\[0\] _04936_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_51_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_16
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12522_ _130_\[20\] _128_\[20\] _06291_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__mux2_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12453_ _132_\[19\] _130_\[19\] _06258_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__mux2_1
X_11404_ _149_\[29\] _132_\[29\] VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__or2_1
X_12384_ _132_\[18\] _134_\[18\] _06219_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__mux2_1
XFILLER_126_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11335_ _05397_ _05398_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__nand2_1
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11266_ _05337_ _05338_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10217_ _04580_ _04584_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__nor2_1
XFILLER_79_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13005_ clknet_leaf_14_clk _00224_ VGND VGND VPWR VPWR _240_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11197_ _05278_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10148_ _03935_ _04085_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__nor2_1
XFILLER_67_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10079_ _03868_ _04454_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__nand2_1
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13907_ clknet_leaf_95_clk _01126_ VGND VGND VPWR VPWR _122_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13838_ clknet_leaf_98_clk _01057_ VGND VGND VPWR VPWR _126_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13769_ clknet_leaf_58_clk _00988_ VGND VGND VPWR VPWR _130_\[9\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_42_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07290_ _01811_ _01834_ _01848_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__nor3_1
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09931_ _04311_ _04312_ _03945_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__a21o_1
XFILLER_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09862_ _04222_ _04225_ _04245_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _03954_ _03876_ _04179_ _01235_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__a211oi_1
XFILLER_133_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08813_ _03233_ _03235_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__xor2_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _228_\[10\] _231_\[10\] _03168_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__o21a_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08675_ _02839_ _02801_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__xnor2_2
XFILLER_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _02170_ _02172_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__nor2_1
XFILLER_54_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07557_ _182_\[14\] _01650_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__or2_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
X_06508_ _190_\[3\] _01220_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__xor2_1
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07488_ _01664_ _01620_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09227_ _02849_ _01426_ _03379_ _03637_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__o211a_1
XFILLER_135_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09158_ _02842_ _01426_ _03379_ _03570_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__o211a_1
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08109_ _234_\[8\] _02564_ _02629_ _02631_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__a211o_1
X_09089_ _03368_ _03501_ _03503_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__o21ai_2
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11120_ net8 _05190_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__and2_1
XFILLER_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11051_ _164_\[21\] _03512_ _04636_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__mux2_1
XFILLER_130_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10002_ _04377_ _04378_ _142_\[20\] VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__a21oi_1
XFILLER_103_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11953_ net13 _05952_ _05852_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__mux2_1
X_11884_ _05864_ _05869_ _05879_ _05889_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__o31a_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10904_ _164_\[3\] _167_\[3\] _05064_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__mux2_1
X_13623_ clknet_leaf_50_clk _00842_ VGND VGND VPWR VPWR _140_\[23\] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_2_3_0_clk clknet_1_1_0_clk VGND VGND VPWR VPWR clknet_2_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10835_ _170_\[15\] _05002_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_24_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
X_13554_ clknet_leaf_74_clk _00773_ VGND VGND VPWR VPWR _149_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10766_ _04971_ _04976_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__or2_1
X_13485_ clknet_leaf_36_clk _00704_ VGND VGND VPWR VPWR _158_\[3\] sky130_fd_sc_hd__dfxtp_1
X_12505_ _130_\[12\] _128_\[12\] _06280_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__mux2_1
X_10697_ _170_\[7\] _173_\[7\] _04830_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__mux2_1
XFILLER_126_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12436_ _132_\[11\] _130_\[11\] _06247_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__mux2_1
XFILLER_113_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12367_ _132_\[10\] _134_\[10\] _06208_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__mux2_1
X_12298_ _06180_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11318_ _05368_ _05373_ _05376_ _05375_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__a31o_1
XFILLER_4_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11249_ _05313_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__nand2_1
XFILLER_113_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06790_ _179_\[5\] _01299_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__or2_1
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08460_ _02890_ _02893_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__xnor2_1
X_07411_ _01949_ _01964_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__nand2_1
XFILLER_63_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08391_ _228_\[20\] _02771_ _02834_ _02837_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__o211a_1
X_07342_ _01897_ _01898_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_15_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07273_ _01830_ _01831_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09012_ _03396_ _03359_ _03395_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__nand3b_1
XFILLER_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09914_ _04195_ _04202_ _04204_ _04267_ _04294_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__a311o_1
XFILLER_59_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09845_ _03896_ _03927_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__nand2_1
XFILLER_113_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _03872_ _04057_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__nand2_1
XFILLER_85_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06988_ _243_\[26\] _01583_ _01557_ _01589_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__a211o_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _03134_ _03135_ _03152_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__and3_1
XFILLER_27_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08658_ _03070_ _03085_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__xor2_2
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _02151_ _02154_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__nand2_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08589_ _03015_ _03018_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10620_ _173_\[14\] _176_\[14\] _01215_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__mux2_1
XFILLER_50_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10551_ _179_\[25\] _04799_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__or2_1
XFILLER_50_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10482_ _173_\[4\] _04735_ _04779_ _04740_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__o211a_1
X_13270_ clknet_leaf_7_clk _00489_ VGND VGND VPWR VPWR _179_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12221_ _138_\[5\] _136_\[5\] _06134_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__mux2_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12152_ _140_\[4\] _138_\[4\] _06101_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__mux2_1
XFILLER_123_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12083_ _06067_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__clkbuf_1
X_11103_ _01254_ _05205_ _05194_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__a21oi_1
XFILLER_123_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11034_ _04855_ _05160_ _05161_ _01436_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__a211o_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12985_ clknet_leaf_14_clk _00204_ VGND VGND VPWR VPWR _243_\[25\] sky130_fd_sc_hd__dfxtp_1
X_11936_ _05924_ _05928_ _05922_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11867_ _140_\[30\] _140_\[0\] VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13606_ clknet_leaf_52_clk _00825_ VGND VGND VPWR VPWR _140_\[6\] sky130_fd_sc_hd__dfxtp_1
X_11798_ _05811_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__clkbuf_1
X_10818_ _167_\[10\] _170_\[10\] _04995_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__mux2_1
XFILLER_32_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13537_ clknet_leaf_66_clk _00756_ VGND VGND VPWR VPWR _149_\[1\] sky130_fd_sc_hd__dfxtp_1
X_10749_ _173_\[22\] _04953_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__or2_1
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13468_ clknet_leaf_122_clk _00687_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dfxtp_4
XFILLER_142_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12419_ _132_\[3\] _130_\[3\] _06201_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__mux2_1
XFILLER_99_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13399_ clknet_leaf_124_clk _00618_ VGND VGND VPWR VPWR _167_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07960_ _02494_ _02495_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__xnor2_1
X_06911_ _01448_ _01534_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__or2_1
XFILLER_68_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07891_ _02385_ _02386_ _02427_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__and3_1
X_09630_ _246_\[5\] _01313_ _03914_ _243_\[5\] _01445_ VGND VGND VPWR VPWR _04023_
+ sky130_fd_sc_hd__o221a_1
X_06842_ _246_\[17\] _01422_ _01481_ _01484_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__o211a_1
XFILLER_56_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09561_ _01282_ _01279_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__or2b_1
X_06773_ _246_\[1\] _01422_ _01425_ _01431_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__o211a_1
XFILLER_83_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08512_ _02932_ _02934_ _02943_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__o21ai_1
X_09492_ _03889_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__clkbuf_4
XFILLER_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08443_ _01719_ _02877_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__nand2_1
XFILLER_51_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08374_ _01411_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07325_ _01881_ _01882_ _01354_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__o21a_1
XFILLER_137_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07256_ _01786_ _01803_ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__o21a_1
XFILLER_105_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07187_ _182_\[2\] _01608_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__nor2_1
XFILLER_105_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09828_ _01242_ _01280_ _04080_ _04087_ _03983_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__a32o_1
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09759_ _04128_ _04147_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _122_\[10\] _120_\[10\] _06423_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__mux2_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _05741_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__clkbuf_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _05678_ _05679_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__nand2_1
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10603_ _176_\[9\] VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__inv_2
X_13322_ clknet_leaf_22_clk _00541_ VGND VGND VPWR VPWR _173_\[4\] sky130_fd_sc_hd__dfxtp_1
X_11583_ _118_\[3\] _05617_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10534_ _176_\[20\] _179_\[20\] _04790_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__mux2_1
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10465_ _176_\[0\] _179_\[0\] _04743_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__mux2_1
X_13253_ clknet_leaf_5_clk _00472_ VGND VGND VPWR VPWR _182_\[31\] sky130_fd_sc_hd__dfxtp_1
X_12204_ _140_\[29\] _138_\[29\] _06123_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__mux2_1
XFILLER_123_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13184_ clknet_leaf_31_clk _00403_ _00105_ VGND VGND VPWR VPWR _195_\[0\] sky130_fd_sc_hd__dfrtp_2
X_10396_ _179_\[12\] _04684_ _04705_ _04717_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__o211a_1
XFILLER_135_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12135_ _140_\[28\] _142_\[28\] _06090_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__mux2_1
XFILLER_97_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12066_ net24 _01274_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__and2_1
XFILLER_49_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11017_ _03125_ _04682_ _04627_ net66 VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_65_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12968_ clknet_leaf_43_clk _00187_ VGND VGND VPWR VPWR _243_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11919_ _140_\[28\] _05920_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__xnor2_1
X_12899_ clknet_leaf_89_clk _00123_ VGND VGND VPWR VPWR _116_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07110_ _01670_ _01682_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__or2_1
X_08090_ _231_\[3\] _02611_ _01695_ _02617_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__o211a_1
X_07041_ _237_\[8\] VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__buf_6
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08992_ _02823_ _02845_ _03379_ _03409_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__o211a_1
X_07943_ _182_\[27\] _01694_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__nor2_1
XFILLER_83_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07874_ _02172_ _02286_ _02407_ _02412_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__o31ai_2
XFILLER_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09613_ _03901_ _04006_ _03873_ _01234_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__a31o_1
X_06825_ _246_\[13\] _01422_ _01425_ _01471_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__o211a_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09544_ _03871_ _03932_ _03940_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__o21ai_1
X_06756_ _392_\[1\] _01415_ net34 VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__a21o_2
XFILLER_43_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09475_ _01280_ _01283_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__nand2b_4
X_06687_ _01375_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08426_ _228_\[28\] _02838_ _02861_ _02864_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__a211o_1
X_08357_ _225_\[13\] VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__clkbuf_4
XFILLER_20_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07308_ _01661_ _01642_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__xnor2_1
X_08288_ _228_\[28\] _02733_ _02723_ _02758_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__o211a_1
XFILLER_137_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07239_ _01520_ _01777_ _01798_ _01799_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__o211a_1
X_10250_ _04437_ _04107_ _04616_ _01233_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__o211a_1
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10181_ _04527_ _04537_ _04550_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__a21oi_1
XFILLER_59_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13940_ clknet_leaf_92_clk _01159_ VGND VGND VPWR VPWR _120_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13871_ clknet_leaf_95_clk _01090_ VGND VGND VPWR VPWR _124_\[15\] sky130_fd_sc_hd__dfxtp_1
X_12822_ _118_\[3\] _120_\[3\] _06451_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__mux2_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12753_ _122_\[2\] _120_\[2\] _06412_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__mux2_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11704_ _05725_ _05726_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__nand2_1
XFILLER_70_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _124_\[1\] _122_\[1\] _06379_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__mux2_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11635_ _05663_ _05664_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__nand2_1
X_11566_ _116_\[15\] _05601_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__nand2_1
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10517_ _176_\[15\] _179_\[15\] _04790_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__mux2_1
X_13305_ clknet_leaf_6_clk _00524_ VGND VGND VPWR VPWR _176_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11497_ _118_\[11\] _05540_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__xnor2_1
X_13236_ clknet_leaf_7_clk _00455_ VGND VGND VPWR VPWR _182_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10448_ _176_\[26\] _04725_ _04755_ _04728_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__a211o_1
X_10379_ _182_\[7\] _04696_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__or2_1
X_13167_ clknet_leaf_108_clk _00386_ VGND VGND VPWR VPWR _225_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12118_ _140_\[20\] _142_\[20\] _06079_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__mux2_1
XFILLER_2_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13098_ clknet_leaf_106_clk _00317_ VGND VGND VPWR VPWR _231_\[10\] sky130_fd_sc_hd__dfxtp_1
X_12049_ _140_\[14\] _140_\[16\] VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__nand2_1
XFILLER_84_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06610_ _392_\[4\] _01206_ _01246_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__or3_4
XFILLER_92_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07590_ _02108_ _02110_ _02107_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06541_ _392_\[1\] _392_\[0\] _01209_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__nand3_2
XFILLER_34_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09260_ _02852_ _03032_ _03309_ _03669_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__a211o_1
XFILLER_33_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08211_ _164_\[6\] _02701_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__or2_1
XFILLER_21_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09191_ _03467_ _03474_ _03542_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__o21bai_1
XFILLER_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08142_ _167_\[18\] _02652_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__or2_1
X_08073_ _182_\[31\] _01707_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07024_ _237_\[4\] VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__buf_4
XFILLER_142_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08975_ _228_\[17\] _231_\[17\] _03392_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__o21a_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07926_ _02462_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__inv_2
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07857_ _02394_ _02395_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__and2_1
X_06808_ _01444_ _01458_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__nand2_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07788_ _185_\[22\] _234_\[22\] VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__nand2_1
X_09527_ _03874_ _01291_ _03923_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__or3_1
X_06739_ net34 VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__inv_2
XFILLER_25_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09458_ _03860_ _03861_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__xnor2_2
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08409_ _228_\[24\] _02838_ _02810_ _02851_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__a211o_1
X_09389_ _03750_ _03753_ _03793_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__and3_1
XFILLER_137_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11420_ _05471_ _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11351_ _05411_ _05412_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__nand2_1
X_10302_ _179_\[12\] _04646_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__or2_1
XFILLER_4_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11282_ _05342_ _05344_ _05350_ _05352_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__a31o_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10233_ _246_\[30\] _01316_ _04409_ _243_\[30\] _01516_ VGND VGND VPWR VPWR _04601_
+ sky130_fd_sc_hd__o221a_2
X_13021_ clknet_leaf_3_clk _00240_ VGND VGND VPWR VPWR _240_\[29\] sky130_fd_sc_hd__dfxtp_1
X_10164_ _185_\[26\] _03867_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__or2_1
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10095_ _04467_ _04468_ _04469_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__a21o_1
XFILLER_75_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13923_ clknet_leaf_70_clk _01142_ VGND VGND VPWR VPWR _120_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13854_ clknet_leaf_69_clk _01073_ VGND VGND VPWR VPWR _126_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12805_ _122_\[27\] _120_\[27\] _01367_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__mux2_1
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13785_ clknet_leaf_76_clk _01004_ VGND VGND VPWR VPWR _130_\[25\] sky130_fd_sc_hd__dfxtp_1
X_10997_ _164_\[31\] _05107_ _04865_ _05139_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__o211a_1
X_12736_ _124_\[26\] _122_\[26\] _06401_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__mux2_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12667_ _126_\[25\] _124_\[25\] _06368_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__mux2_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11618_ _05639_ _05648_ _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__or3_1
XFILLER_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12598_ _128_\[24\] _126_\[24\] _06335_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__mux2_1
XFILLER_51_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11549_ _05578_ _05580_ _05576_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__o21ai_1
XFILLER_116_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13219_ clknet_leaf_41_clk _00438_ VGND VGND VPWR VPWR _185_\[29\] sky130_fd_sc_hd__dfxtp_2
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _02404_ _03184_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__nand2_1
X_07711_ _02213_ _02239_ _02253_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__nor3_1
X_08691_ _03100_ _03117_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07642_ _02184_ _02187_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__xor2_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07573_ _02117_ _02120_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__or2_1
X_09312_ _03718_ _03719_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__and2_1
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06524_ _01232_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__clkbuf_4
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09243_ _03651_ _03652_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__or2_1
XFILLER_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09174_ _03583_ _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__xor2_1
XFILLER_135_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08125_ _231_\[13\] _02611_ _02641_ _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__o211a_1
XFILLER_107_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08056_ _02586_ _02588_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07007_ _01568_ _01602_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__or2_1
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput38 net38 VGND VGND VPWR VPWR dout[11] sky130_fd_sc_hd__buf_2
Xoutput49 net49 VGND VGND VPWR VPWR dout[21] sky130_fd_sc_hd__buf_2
XFILLER_143_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08958_ _02404_ _03376_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__nand2_1
XFILLER_57_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07909_ _01355_ _02439_ _02440_ _02446_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__a31o_1
X_08889_ _01417_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__buf_6
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10920_ net65 _05068_ _05085_ _05086_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__a211o_1
XFILLER_112_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10851_ _167_\[19\] _05022_ _05009_ _05037_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__o211a_1
X_13570_ clknet_leaf_34_clk _00789_ VGND VGND VPWR VPWR _142_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10782_ _167_\[31\] _04986_ _04988_ _04952_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__a211o_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12521_ _06297_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__clkbuf_1
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12452_ _06261_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__clkbuf_1
X_11403_ _149_\[29\] _132_\[29\] VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__nand2_1
XFILLER_138_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12383_ _06225_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__clkbuf_1
X_11334_ _05381_ _05386_ _05389_ _05388_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__a31o_1
XFILLER_4_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11265_ _05328_ _05331_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__nand2_1
XFILLER_4_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10216_ _04580_ _04584_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__and2_1
X_13004_ clknet_leaf_17_clk _00223_ VGND VGND VPWR VPWR _240_\[12\] sky130_fd_sc_hd__dfxtp_1
X_11196_ _152_\[2\] _05277_ _01362_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__mux2_1
XFILLER_95_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10147_ _01232_ _04333_ _04366_ _04518_ _04362_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__o32a_1
XFILLER_121_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10078_ _04449_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13906_ clknet_leaf_96_clk _01125_ VGND VGND VPWR VPWR _122_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13837_ clknet_leaf_95_clk _01056_ VGND VGND VPWR VPWR _126_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13768_ clknet_leaf_58_clk _00987_ VGND VGND VPWR VPWR _130_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_12719_ _01392_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__buf_4
XFILLER_31_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13699_ clknet_leaf_59_clk _00918_ VGND VGND VPWR VPWR _134_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09930_ _04295_ _04296_ _04310_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__nand3_1
XFILLER_131_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09861_ _04222_ _04225_ _04245_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__and3_1
XFILLER_124_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _03934_ _03923_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__nor2_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08812_ _03198_ _03200_ _03234_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__o21ai_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _228_\[10\] _231_\[10\] _02801_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__a21o_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08674_ _01930_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__clkinv_2
XFILLER_66_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _02108_ _02110_ _02135_ _02136_ _02171_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__o311a_1
XFILLER_53_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07556_ _02101_ _02104_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__xor2_1
XFILLER_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06507_ _190_\[2\] _190_\[1\] _190_\[0\] _01213_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__and4_1
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07487_ _02037_ _02012_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__or2_1
XFILLER_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09226_ _01428_ _03607_ _03636_ _01495_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__a211o_1
XFILLER_10_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09157_ _01421_ _03569_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__nand2_1
X_08108_ _231_\[8\] _02611_ _01695_ _02630_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__o211a_1
X_09088_ _03426_ _03457_ _03458_ _03502_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__o211a_1
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08039_ _01632_ _01616_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__xnor2_2
XFILLER_131_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11050_ _03478_ _04855_ _04628_ net48 _05171_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__o221a_1
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10001_ _142_\[20\] _04377_ _04378_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__and3_1
XFILLER_89_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11952_ _05946_ _05951_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__xor2_1
XFILLER_45_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11883_ _05867_ _05876_ _05877_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__a21o_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10903_ net58 _05068_ _05074_ _05035_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__a211o_1
X_13622_ clknet_leaf_49_clk _00841_ VGND VGND VPWR VPWR _140_\[22\] sky130_fd_sc_hd__dfxtp_2
X_10834_ _04682_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__buf_2
X_13553_ clknet_leaf_79_clk _00772_ VGND VGND VPWR VPWR _149_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12504_ _06288_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10765_ _170_\[27\] _173_\[27\] _04936_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__mux2_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13484_ clknet_leaf_36_clk _00703_ VGND VGND VPWR VPWR _158_\[2\] sky130_fd_sc_hd__dfxtp_1
X_10696_ _167_\[6\] _04925_ _04927_ _04891_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__o211a_1
XFILLER_138_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12435_ _06252_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12366_ _06216_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11317_ _05381_ _05382_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__nand2_1
X_12297_ _136_\[9\] _134_\[9\] _06178_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__mux2_1
XFILLER_113_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11248_ _05314_ _05316_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__or2_1
X_11179_ _01361_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__clkbuf_4
XFILLER_95_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07410_ _01962_ _01963_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__and2_1
X_08390_ _02002_ _02836_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__or2_1
XFILLER_23_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07341_ _185_\[7\] _234_\[7\] VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__or2_1
X_07272_ _01822_ _01823_ _01821_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__o21a_1
XFILLER_145_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09011_ _03426_ _03427_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__and2_1
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09913_ _04290_ _04287_ _04294_ _04269_ _04288_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__o221a_1
X_09844_ _142_\[13\] _04228_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _04010_ _03936_ _04002_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__o21a_1
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06987_ _240_\[26\] _01565_ _01558_ _01588_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__o211a_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08726_ _03136_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__xor2_1
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08657_ _03081_ _03084_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__xnor2_2
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _02151_ _02154_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__or2_1
X_08588_ _03016_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__nor2_1
XFILLER_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07539_ _01671_ _01626_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__xnor2_1
X_10550_ _173_\[24\] _04774_ _04827_ _04777_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__a211o_1
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10481_ _04766_ _04778_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__or2_1
X_09209_ _03618_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__nand2_1
X_12220_ _06139_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12151_ _06103_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12082_ _140_\[3\] _142_\[3\] _06005_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__mux2_1
X_11102_ _05203_ _158_\[3\] VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__or2b_1
XFILLER_123_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11033_ _03306_ _04631_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__nor2_1
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12984_ clknet_leaf_14_clk _00203_ VGND VGND VPWR VPWR _243_\[24\] sky130_fd_sc_hd__dfxtp_1
X_11935_ _05934_ _05935_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__nand2_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13605_ clknet_leaf_53_clk _00824_ VGND VGND VPWR VPWR _140_\[5\] sky130_fd_sc_hd__dfxtp_1
X_11866_ _05873_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__clkbuf_1
X_11797_ _142_\[6\] _05810_ _05765_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__mux2_1
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10817_ _164_\[9\] _04986_ _05013_ _05001_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__a211o_1
X_13536_ clknet_leaf_68_clk _00755_ VGND VGND VPWR VPWR _149_\[0\] sky130_fd_sc_hd__dfxtp_1
X_10748_ _167_\[21\] _04925_ _04964_ _04939_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__o211a_1
XFILLER_9_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13467_ clknet_leaf_128_clk _00686_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dfxtp_2
XFILLER_145_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12418_ _06243_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__clkbuf_1
X_10679_ _170_\[2\] _173_\[2\] _04830_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__mux2_1
XFILLER_138_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13398_ clknet_leaf_125_clk _00617_ VGND VGND VPWR VPWR _167_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12349_ _06207_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06910_ _176_\[4\] _240_\[4\] _01449_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__mux2_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07890_ _02385_ _02386_ _02427_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__a21oi_1
X_06841_ _01444_ _01483_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__nand2_1
XFILLER_68_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09560_ _01234_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__nand2_1
X_06772_ _01426_ _01430_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__nand2_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09491_ _195_\[2\] _195_\[1\] VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__or2_1
XFILLER_82_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08511_ _170_\[2\] _02776_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__nand2_1
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08442_ _01714_ _02876_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08373_ _225_\[17\] VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__clkbuf_4
X_07324_ _01864_ _01880_ _01879_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__a21oi_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07255_ _01813_ _01814_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07186_ _01747_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__inv_2
XFILLER_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_2_0_clk clknet_1_1_0_clk VGND VGND VPWR VPWR clknet_2_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_59_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09827_ _03898_ _03880_ _04132_ _03888_ _01236_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__a221o_1
XFILLER_101_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09758_ _04144_ _04146_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__nand2_1
XFILLER_86_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08709_ _03100_ _03117_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__or2b_1
X_09689_ _03896_ _03888_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__nand2_2
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _149_\[31\] _05740_ _05625_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__mux2_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _116_\[24\] _05677_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__or2_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10602_ _04861_ _04862_ _04863_ _04823_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__o211a_1
X_11582_ _118_\[20\] _118_\[24\] VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13321_ clknet_leaf_18_clk _00540_ VGND VGND VPWR VPWR _173_\[3\] sky130_fd_sc_hd__dfxtp_2
X_10533_ _173_\[19\] _04780_ _04815_ _04785_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__o211a_1
XFILLER_10_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10464_ _04681_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__buf_2
X_13252_ clknet_leaf_5_clk _00471_ VGND VGND VPWR VPWR _182_\[30\] sky130_fd_sc_hd__dfxtp_1
X_12203_ _06130_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__clkbuf_1
X_10395_ _182_\[12\] _04696_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__or2_1
X_13183_ clknet_leaf_120_clk _00402_ VGND VGND VPWR VPWR _225_\[31\] sky130_fd_sc_hd__dfxtp_1
X_12134_ _06094_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12065_ _06038_ _06052_ _06042_ _06051_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__a211o_1
XFILLER_49_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11016_ net65 _04629_ _05150_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__o21a_1
XFILLER_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12967_ clknet_leaf_17_clk _00186_ VGND VGND VPWR VPWR _243_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11918_ _140_\[3\] _140_\[5\] VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__xnor2_1
X_12898_ clknet_leaf_73_clk _00122_ VGND VGND VPWR VPWR _116_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11849_ _152_\[11\] _05856_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__or2_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13519_ clknet_leaf_78_clk _00738_ VGND VGND VPWR VPWR _152_\[15\] sky130_fd_sc_hd__dfxtp_1
X_07040_ _240_\[7\] _01583_ _01607_ _01628_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__a211o_1
XFILLER_114_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08991_ _01520_ _03402_ _03408_ _02355_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__a211o_1
XFILLER_141_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07942_ _01690_ _02448_ _02419_ _02478_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__o211a_1
X_07873_ _182_\[23\] _01681_ _02411_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__a21oi_1
X_09612_ _01241_ _04005_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__nor2_2
X_06824_ _01444_ _01470_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__nand2_1
XFILLER_96_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09543_ _03933_ _03934_ _03937_ _03939_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__a31o_1
XFILLER_95_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06755_ _392_\[0\] _01210_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__nor2_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09474_ _01234_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__buf_2
X_06686_ _118_\[8\] _116_\[8\] _01370_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__mux2_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08425_ _02862_ _01801_ _02824_ _02863_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__o211a_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08356_ _02711_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__clkbuf_4
X_07307_ _01846_ _01847_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__and2b_1
X_08287_ _164_\[28\] _02736_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__or2_1
XFILLER_118_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07238_ _01412_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__buf_4
XFILLER_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07169_ _01714_ _01716_ _01715_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__a21boi_1
XFILLER_133_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10180_ _04527_ _04537_ _04550_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__and3_1
XFILLER_105_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13870_ clknet_leaf_98_clk _01089_ VGND VGND VPWR VPWR _124_\[14\] sky130_fd_sc_hd__dfxtp_1
X_12821_ _06454_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12752_ _06418_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__clkbuf_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12683_ _06382_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__clkbuf_1
X_11703_ _116_\[29\] _05722_ _05723_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__nand3_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11634_ _116_\[22\] _05662_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__or2_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11565_ _116_\[15\] _05601_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__nor2_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11496_ _118_\[26\] _118_\[15\] VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__xnor2_1
X_10516_ _173_\[14\] _04774_ _04803_ _04777_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__a211o_1
X_13304_ clknet_leaf_9_clk _00523_ VGND VGND VPWR VPWR _176_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13235_ clknet_leaf_25_clk _00454_ VGND VGND VPWR VPWR _182_\[13\] sky130_fd_sc_hd__dfxtp_1
X_10447_ _179_\[26\] _04721_ _04751_ _04754_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__o211a_1
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10378_ _04685_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__clkbuf_4
X_13166_ clknet_leaf_106_clk _00385_ VGND VGND VPWR VPWR _225_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12117_ _06085_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13097_ clknet_leaf_116_clk _00316_ VGND VGND VPWR VPWR _231_\[9\] sky130_fd_sc_hd__dfxtp_1
X_12048_ _140_\[14\] _140_\[16\] VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__or2_1
XFILLER_78_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06540_ _392_\[4\] _01246_ _01248_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08210_ _231_\[5\] _02690_ _02664_ _02703_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__a211o_1
XFILLER_21_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09190_ _03469_ _03510_ _03541_ _03593_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__or4bb_1
X_08141_ _234_\[17\] _02646_ _02629_ _02654_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__a211o_1
X_08072_ _02557_ _02567_ _02568_ _02565_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__o31a_1
X_07023_ _01405_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__clkbuf_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08974_ _228_\[17\] _231_\[17\] _02823_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__a21o_1
X_07925_ _02428_ _02449_ _02461_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__o21a_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07856_ _02368_ _02381_ _02393_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__or3_1
X_06807_ _243_\[9\] _01428_ _01457_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07787_ _185_\[22\] _234_\[22\] VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__or2_1
X_09526_ _195_\[1\] _195_\[0\] VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__nor2_1
X_06738_ net34 VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__inv_2
X_09457_ _170_\[31\] _02871_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06669_ _01364_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08408_ _02849_ _01801_ _02824_ _02850_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__o211a_1
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09388_ _03750_ _03753_ _03793_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08339_ _225_\[9\] VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__clkbuf_4
XFILLER_137_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11350_ _05395_ _05400_ _05403_ _05402_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__a31o_1
XFILLER_137_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10301_ _179_\[11\] _04629_ _04655_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__a21o_1
XFILLER_4_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11281_ _01367_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__buf_4
XFILLER_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13020_ clknet_leaf_13_clk _00239_ VGND VGND VPWR VPWR _240_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10232_ _01233_ _04595_ _04596_ _04599_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__o31a_1
XFILLER_105_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10163_ _04529_ _04534_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__xor2_1
X_10094_ _04467_ _04468_ _03867_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__o21ai_1
X_13922_ clknet_leaf_70_clk _01141_ VGND VGND VPWR VPWR _120_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13853_ clknet_leaf_72_clk _01072_ VGND VGND VPWR VPWR _126_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12804_ _06445_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__clkbuf_1
X_13784_ clknet_leaf_76_clk _01003_ VGND VGND VPWR VPWR _130_\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10996_ _167_\[31\] _04867_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__or2_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _06409_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12666_ _06373_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__clkbuf_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11617_ _05631_ _05633_ _05638_ _05629_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__o211a_1
XFILLER_30_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12597_ _06337_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11548_ _05585_ _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__or2b_1
XFILLER_11_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11479_ _149_\[6\] _05524_ _05439_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__mux2_1
XFILLER_124_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13218_ clknet_leaf_38_clk _00437_ VGND VGND VPWR VPWR _185_\[28\] sky130_fd_sc_hd__dfxtp_4
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13149_ clknet_leaf_119_clk _00368_ VGND VGND VPWR VPWR _228_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _02213_ _02239_ _02253_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__o21a_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08690_ _03115_ _03116_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07641_ _02185_ _02186_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__nand2_1
XFILLER_81_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07572_ _02118_ _02119_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__nand2_1
XFILLER_19_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06523_ _01231_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__buf_2
XFILLER_80_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09311_ _03709_ _03711_ _03717_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__nand3_1
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09242_ _03615_ _03619_ _03650_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__and3_1
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09173_ _228_\[23\] _231_\[23\] _03584_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__o21ai_2
X_08124_ _167_\[13\] _02616_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__or2_1
XFILLER_119_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08055_ _02518_ _02523_ _02552_ _02553_ _02587_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__o41a_1
XFILLER_89_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07006_ _173_\[0\] _237_\[0\] _01569_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__mux2_1
Xoutput39 net39 VGND VGND VPWR VPWR dout[12] sky130_fd_sc_hd__buf_2
XFILLER_89_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08957_ _03372_ _03375_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__xnor2_2
XFILLER_29_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07908_ _01778_ _02445_ _01412_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__o21ai_2
X_08888_ _02814_ _03032_ _02861_ _03308_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__a211o_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07839_ _01856_ _02359_ _02378_ _02355_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__a211o_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10850_ _170_\[19\] _05036_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__or2_1
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09509_ _01240_ _01280_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__or2_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10781_ _170_\[31\] _04980_ _04958_ _04987_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__o211a_1
XFILLER_24_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _130_\[19\] _128_\[19\] _06291_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__mux2_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12451_ _132_\[18\] _130_\[18\] _06258_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__mux2_1
XFILLER_138_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11402_ _05457_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12382_ _132_\[17\] _134_\[17\] _06219_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__mux2_1
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11333_ _05396_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__inv_2
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11264_ _05335_ _05336_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__or2b_1
X_10215_ _04582_ _04583_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__nor2_1
XFILLER_106_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13003_ clknet_leaf_14_clk _00222_ VGND VGND VPWR VPWR _240_\[11\] sky130_fd_sc_hd__dfxtp_1
X_11195_ _05273_ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10146_ _04027_ _03976_ _04103_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__o21a_1
XFILLER_67_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10077_ _04451_ _04452_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__or2_1
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13905_ clknet_leaf_95_clk _01124_ VGND VGND VPWR VPWR _122_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13836_ clknet_leaf_98_clk _01055_ VGND VGND VPWR VPWR _126_\[12\] sky130_fd_sc_hd__dfxtp_1
X_13767_ clknet_leaf_60_clk _00986_ VGND VGND VPWR VPWR _130_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10979_ _164_\[25\] _05107_ _05094_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__o211a_1
XFILLER_16_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12718_ _06400_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__clkbuf_1
X_13698_ clknet_leaf_59_clk _00917_ VGND VGND VPWR VPWR _134_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12649_ _06364_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09860_ _04243_ _04244_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__and2b_1
XFILLER_140_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _04002_ _01292_ _04027_ _04177_ _01235_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__o311a_1
XFILLER_98_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08811_ _03201_ _03203_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__or2b_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08742_ _03164_ _03166_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__xnor2_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08673_ _03095_ _03099_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__and2_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07624_ _02135_ _01650_ _182_\[14\] VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__nand3b_1
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07555_ _02035_ _02052_ _02078_ _02103_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__a31o_1
XFILLER_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06506_ _190_\[2\] _190_\[1\] _190_\[0\] _190_\[3\] VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__or4b_1
X_07486_ _02009_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__inv_2
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09225_ _03628_ _03634_ _03635_ _01523_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__o211a_1
XFILLER_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09156_ _03544_ _03568_ _01354_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__mux2_1
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_110_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_110_clk sky130_fd_sc_hd__clkbuf_16
X_08107_ _167_\[8\] _02616_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__or2_1
X_09087_ _03500_ _03430_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__or2b_1
XFILLER_135_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08038_ _02548_ _02549_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__and2b_1
XFILLER_116_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10000_ _246_\[20\] _01315_ _01301_ _179_\[20\] VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__o22a_1
XFILLER_107_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09989_ _04361_ _04362_ _04364_ _04255_ _04367_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__o221a_1
XFILLER_76_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11951_ _05909_ _05948_ _05950_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__o21a_1
XFILLER_29_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11882_ _05886_ _05887_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__nand2_1
XFILLER_83_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10902_ _164_\[2\] _05059_ _05043_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__o211a_1
X_13621_ clknet_leaf_49_clk _00840_ VGND VGND VPWR VPWR _140_\[21\] sky130_fd_sc_hd__dfxtp_2
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10833_ _164_\[14\] _04986_ _05024_ _05001_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__a211o_1
XFILLER_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13552_ clknet_leaf_84_clk _00771_ VGND VGND VPWR VPWR _149_\[16\] sky130_fd_sc_hd__dfxtp_1
X_10764_ _167_\[26\] _04945_ _04975_ _04952_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__a211o_1
X_12503_ _130_\[11\] _128_\[11\] _06280_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__mux2_1
XFILLER_40_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13483_ clknet_leaf_35_clk _00702_ VGND VGND VPWR VPWR _158_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10695_ _04888_ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__or2_1
XFILLER_145_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12434_ _132_\[10\] _130_\[10\] _06247_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__mux2_1
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12365_ _132_\[9\] _134_\[9\] _06208_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__mux2_1
XFILLER_66_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_101_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_101_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_126_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11316_ _149_\[18\] _132_\[18\] VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__or2_1
XFILLER_5_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12296_ _06179_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11247_ _05320_ _05321_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__or2b_1
XFILLER_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11178_ _01368_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__clkbuf_4
X_10129_ _04501_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__inv_2
XFILLER_95_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13819_ clknet_leaf_71_clk _01038_ VGND VGND VPWR VPWR _128_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07340_ _185_\[7\] _234_\[7\] VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__nand2_1
XFILLER_16_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07271_ _01828_ _01829_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__nand2_1
X_09010_ _03410_ _03411_ _03425_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__or3_1
XFILLER_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09912_ _04266_ _04289_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__or2_1
XFILLER_113_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09843_ _246_\[13\] _01315_ _04129_ _243_\[13\] _01469_ VGND VGND VPWR VPWR _04228_
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _04051_ _04132_ _04160_ _03903_ _04161_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__a221o_1
XFILLER_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06986_ _176_\[26\] _01580_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__or2_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ _03147_ _03150_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__xnor2_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _03082_ _03083_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__nor2_1
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _02152_ _02153_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__nand2_1
X_08587_ _228_\[5\] _231_\[5\] _02784_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__a21oi_2
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07538_ _01645_ _01973_ _01886_ _02087_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__o211a_1
XFILLER_41_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07469_ _02019_ _02020_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__or2b_1
XFILLER_22_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10480_ _176_\[4\] _179_\[4\] _04743_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__mux2_1
X_09208_ _02392_ _03617_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__nand2_1
X_09139_ _03550_ _03551_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__nand2_1
X_12150_ _140_\[3\] _138_\[3\] _06101_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__mux2_1
XFILLER_118_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11101_ net3 _05202_ _05191_ _05203_ _05204_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__a221o_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12081_ _06066_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11032_ net41 _164_\[14\] _01215_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__mux2_1
XFILLER_89_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12983_ clknet_leaf_10_clk _00202_ VGND VGND VPWR VPWR _243_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11934_ _152_\[19\] _05933_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__or2_1
XFILLER_73_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13604_ clknet_leaf_52_clk _00823_ VGND VGND VPWR VPWR _140_\[4\] sky130_fd_sc_hd__dfxtp_2
X_11865_ _142_\[12\] _05872_ _05765_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__mux2_1
XFILLER_26_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11796_ net29 _05776_ _05807_ _05809_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__a22o_1
XFILLER_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10816_ _167_\[9\] _04980_ _05009_ _05012_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__o211a_1
X_13535_ clknet_leaf_66_clk _00754_ VGND VGND VPWR VPWR _152_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10747_ _04888_ _04963_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__or2_1
XFILLER_139_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10678_ _167_\[1\] _04836_ _04913_ _04914_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__a211o_1
X_13466_ clknet_leaf_123_clk _00685_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dfxtp_2
X_12417_ _132_\[2\] _130_\[2\] _06201_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__mux2_1
XFILLER_126_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13397_ clknet_leaf_124_clk _00616_ VGND VGND VPWR VPWR _167_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12348_ _132_\[1\] _134_\[1\] _06090_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__mux2_1
X_12279_ _06170_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06840_ _243_\[17\] _01438_ _01482_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__o21ai_1
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06771_ _243_\[1\] _01428_ _01429_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__o21ai_1
X_09490_ _01282_ _01278_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__nand2b_4
X_08510_ _02940_ _02941_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__nand2_1
XFILLER_91_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08441_ _185_\[0\] _02875_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08372_ _228_\[16\] _02775_ _02810_ _02822_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__a211o_1
X_07323_ _01864_ _01879_ _01880_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__and3_1
X_07254_ _243_\[4\] _240_\[4\] _01616_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__mux2_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07185_ _182_\[2\] _01608_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__nand2_1
XFILLER_145_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09826_ _01236_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__nand2_1
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09757_ _04145_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__inv_2
XFILLER_104_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06969_ _176_\[21\] _240_\[21\] _01569_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__mux2_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08708_ _03116_ _03115_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__or2b_1
XFILLER_27_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09688_ _04075_ _03954_ _03928_ _04077_ _04078_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__a311o_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08639_ _03025_ _03054_ _03058_ _03066_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__a31o_1
XFILLER_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _116_\[24\] _05677_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__nand2_1
X_10601_ _01922_ _04724_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__nand2_1
X_11581_ _05616_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13320_ clknet_leaf_18_clk _00539_ VGND VGND VPWR VPWR _173_\[2\] sky130_fd_sc_hd__dfxtp_2
X_10532_ _04809_ _04814_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__or2_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10463_ _176_\[31\] _04735_ _04765_ _04740_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__o211a_1
X_13251_ clknet_leaf_5_clk _00470_ VGND VGND VPWR VPWR _182_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12202_ _140_\[28\] _138_\[28\] _06123_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__mux2_1
X_10394_ _176_\[11\] _04683_ _04716_ _01419_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__a211o_1
X_13182_ clknet_leaf_103_clk _00401_ VGND VGND VPWR VPWR _225_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12133_ _140_\[27\] _142_\[27\] _06090_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__mux2_1
XFILLER_89_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12064_ _06051_ _06053_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__nand2_1
XFILLER_97_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11015_ _164_\[7\] _04678_ _03069_ _04686_ _04648_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__o221a_1
XFILLER_77_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12966_ clknet_leaf_20_clk _00185_ VGND VGND VPWR VPWR _243_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11917_ _05919_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__clkbuf_1
X_12897_ clknet_leaf_73_clk _00121_ VGND VGND VPWR VPWR _116_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11848_ _152_\[11\] _05856_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__and2_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11779_ _05793_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__inv_2
X_13518_ clknet_leaf_81_clk _00737_ VGND VGND VPWR VPWR _152_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13449_ clknet_leaf_1_clk _00668_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfxtp_2
XFILLER_127_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08990_ _01778_ _03407_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__nor2_1
XFILLER_142_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07941_ _01355_ _02469_ _02470_ _02477_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__a31o_1
X_07872_ _182_\[23\] _01681_ _02349_ _02409_ _02410_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__o221a_1
X_09611_ _04004_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__buf_2
X_06823_ _243_\[13\] _01428_ _01469_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09542_ _01234_ _03903_ _03938_ _03910_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__a31o_1
X_06754_ _243_\[0\] _01409_ _01412_ _01413_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__o211a_1
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09473_ _01230_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__clkbuf_4
X_06685_ _01374_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_90_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_36_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08424_ net56 _01519_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__or2_1
X_08355_ _228_\[12\] _02771_ _02765_ _02809_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__o211a_1
X_07306_ _01811_ _01834_ _01848_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__or3_1
X_08286_ _231_\[27\] _02730_ _02753_ _02757_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__a211o_1
X_07237_ _01778_ _01797_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__nand2_1
XFILLER_20_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07168_ _01727_ _01730_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07099_ _240_\[20\] _01660_ _01653_ _01674_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__o211a_1
XFILLER_133_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09809_ _04194_ _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__nand2_1
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12820_ _118_\[2\] _120_\[2\] _06451_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__mux2_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12751_ _122_\[1\] _120_\[1\] _06412_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__mux2_1
XFILLER_70_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12682_ _124_\[0\] _122_\[0\] _06379_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__mux2_1
XFILLER_91_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_81_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_16
X_11702_ _05724_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__inv_2
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11633_ _116_\[22\] _05662_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__nand2_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11564_ _118_\[18\] _05600_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11495_ _05501_ _05536_ _05537_ _05538_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__o211a_1
X_10515_ _176_\[14\] _04771_ _04751_ _04802_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__o211a_1
X_13303_ clknet_leaf_7_clk _00522_ VGND VGND VPWR VPWR _176_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13234_ clknet_leaf_26_clk _00453_ VGND VGND VPWR VPWR _182_\[12\] sky130_fd_sc_hd__dfxtp_1
X_10446_ _182_\[26\] _04746_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__or2_1
XFILLER_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10377_ _176_\[6\] _04691_ _04704_ _04677_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__o211a_1
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13165_ clknet_leaf_109_clk _00384_ VGND VGND VPWR VPWR _225_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12116_ _140_\[19\] _142_\[19\] _06079_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__mux2_1
X_13096_ clknet_leaf_109_clk _00315_ VGND VGND VPWR VPWR _231_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12047_ _06030_ _06034_ _06032_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__a21oi_1
XFILLER_93_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12949_ clknet_leaf_29_clk _00168_ VGND VGND VPWR VPWR _246_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_72_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_2_1_0_clk clknet_1_0_0_clk VGND VGND VPWR VPWR clknet_2_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_61_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08140_ _231_\[17\] _02649_ _02641_ _02653_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__o211a_1
X_08071_ _02592_ _02602_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07022_ _240_\[3\] _01583_ _01607_ _01614_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__a211o_1
XFILLER_142_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08973_ _03389_ _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07924_ _02459_ _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07855_ _02368_ _02381_ _02393_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__o21ai_1
X_06806_ _179_\[9\] _01300_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__or2_1
XFILLER_83_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07786_ _02326_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__inv_2
XFILLER_37_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09525_ _142_\[1\] _03921_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__xor2_1
XFILLER_83_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06737_ _01402_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_63_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_16
X_06668_ _116_\[1\] _118_\[1\] _01362_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__mux2_1
X_09456_ _03838_ _03840_ _03837_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__a21bo_1
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08407_ net52 _01519_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__or2_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06599_ _01301_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__buf_4
XFILLER_101_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09387_ _03791_ _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__nand2_1
XFILLER_12_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08338_ _228_\[8\] _02771_ _02765_ _02796_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__o211a_1
XFILLER_138_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08269_ _164_\[23\] _228_\[23\] _02687_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__mux2_1
X_10300_ _182_\[11\] _04654_ _04642_ _04650_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__a31o_1
X_11280_ _05342_ _05344_ _05350_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__a21oi_1
X_10231_ _04210_ _04597_ _04598_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__or3_1
XFILLER_118_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10162_ _04531_ _04533_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__nand2_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10093_ _04449_ _04453_ _04447_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__a21boi_1
XFILLER_105_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13921_ clknet_leaf_70_clk _01140_ VGND VGND VPWR VPWR _120_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13852_ clknet_leaf_71_clk _01071_ VGND VGND VPWR VPWR _126_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12803_ _122_\[26\] _120_\[26\] _01367_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__mux2_1
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13783_ clknet_leaf_94_clk _01002_ VGND VGND VPWR VPWR _130_\[23\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_54_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _124_\[25\] _122_\[25\] _06401_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__mux2_1
XFILLER_43_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10995_ net59 _04853_ _05138_ _05117_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__o211a_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12665_ _126_\[24\] _124_\[24\] _06368_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__mux2_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11616_ _05646_ _05647_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__nand2_1
X_12596_ _128_\[23\] _126_\[23\] _06335_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__mux2_1
X_11547_ _116_\[13\] _05584_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__nand2_1
XFILLER_144_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11478_ _05519_ _05523_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13217_ clknet_leaf_38_clk _00436_ VGND VGND VPWR VPWR _185_\[27\] sky130_fd_sc_hd__dfxtp_4
X_10429_ _04712_ _04741_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__or2_1
XFILLER_98_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13148_ clknet_leaf_119_clk _00367_ VGND VGND VPWR VPWR _228_\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13079_ clknet_leaf_100_clk _00298_ VGND VGND VPWR VPWR _234_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07640_ _185_\[17\] _234_\[17\] VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__nand2_1
XFILLER_66_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07571_ _185_\[15\] _234_\[15\] VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__nand2_1
X_06522_ _01230_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_45_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09310_ _03709_ _03711_ _03717_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__a21o_1
XFILLER_80_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09241_ _03615_ _03619_ _03650_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09172_ _228_\[23\] _231_\[23\] _02846_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__a21o_1
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08123_ _01420_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__clkbuf_4
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08054_ _02516_ _02552_ _02553_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__o21bai_1
XFILLER_134_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07005_ _01421_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08956_ _03335_ _03373_ _03374_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__nor3_4
XFILLER_69_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07907_ _02443_ _02444_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__xnor2_2
XFILLER_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08887_ _02380_ _03300_ _03307_ _01439_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__o211a_1
XFILLER_84_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07838_ _02375_ _02376_ _02377_ _01523_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__o211a_1
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09508_ _03904_ _03905_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_36_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_112_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07769_ _243_\[21\] _240_\[21\] _01675_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__mux2_4
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10780_ _173_\[31\] _04953_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__or2_1
XFILLER_80_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09439_ _02868_ _01884_ _03309_ _03843_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__a211o_1
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12450_ _06260_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__clkbuf_1
X_11401_ _152_\[28\] _05456_ _05439_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__mux2_1
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_80 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12381_ _06224_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11332_ _05394_ _05395_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__and2_1
XFILLER_4_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11263_ _149_\[11\] _132_\[11\] VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__nand2_1
XFILLER_137_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11194_ _05274_ _05275_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__and2b_1
X_10214_ _142_\[29\] _04581_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__nor2_1
X_13002_ clknet_leaf_19_clk _00221_ VGND VGND VPWR VPWR _240_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10145_ _04515_ _04516_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__or2_1
XFILLER_79_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10076_ _04393_ _04425_ _04426_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__o21a_1
XFILLER_75_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13904_ clknet_leaf_96_clk _01123_ VGND VGND VPWR VPWR _122_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13835_ clknet_leaf_93_clk _01054_ VGND VGND VPWR VPWR _126_\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_27_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_90_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13766_ clknet_leaf_60_clk _00985_ VGND VGND VPWR VPWR _130_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10978_ _167_\[25\] _04867_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__or2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13697_ clknet_leaf_59_clk _00916_ VGND VGND VPWR VPWR _134_\[1\] sky130_fd_sc_hd__dfxtp_1
X_12717_ _124_\[17\] _122_\[17\] _06390_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__mux2_1
X_12648_ _126_\[16\] _124_\[16\] _06357_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__mux2_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12579_ _128_\[15\] _126_\[15\] _06324_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__mux2_1
XFILLER_117_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08810_ _03230_ _03232_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__xnor2_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _01283_ _03952_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__nand2_1
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08741_ _01960_ _03143_ _03165_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08672_ _03087_ _03096_ _03097_ _03051_ _03098_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__o221a_1
X_07623_ _02168_ _02169_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__or2_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
X_07554_ _02077_ _02102_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__and2_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07485_ _02016_ _02017_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__and2b_1
X_06505_ _01217_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__buf_6
X_09224_ _03628_ _03634_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__nand2_1
XFILLER_22_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09155_ _03564_ _03567_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08106_ _01435_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__clkbuf_4
X_09086_ _03429_ _03500_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__or2_1
XFILLER_135_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08037_ _02567_ _02569_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__xnor2_2
XFILLER_122_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09988_ _01231_ _01236_ _04365_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__or4_1
XFILLER_107_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08939_ _03324_ _03327_ _03323_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__a21oi_2
X_11950_ _05922_ _05949_ _05947_ _05927_ _05934_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__o221a_1
XFILLER_83_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10901_ _167_\[2\] _05036_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__or2_1
X_11881_ _152_\[14\] _05885_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__or2_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13620_ clknet_leaf_46_clk _00839_ VGND VGND VPWR VPWR _140_\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_72_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10832_ _167_\[14\] _05022_ _05009_ _05023_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__o211a_1
X_13551_ clknet_leaf_87_clk _00770_ VGND VGND VPWR VPWR _149_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10763_ _170_\[26\] _04942_ _04958_ _04974_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__o211a_1
XFILLER_13_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12502_ _06287_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13482_ clknet_leaf_35_clk _00701_ VGND VGND VPWR VPWR _158_\[0\] sky130_fd_sc_hd__dfxtp_1
X_10694_ _170_\[6\] _173_\[6\] _04830_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__mux2_1
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12433_ _06251_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__clkbuf_1
X_12364_ _06215_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11315_ _149_\[18\] _132_\[18\] VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__nand2_1
XFILLER_141_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12295_ _136_\[8\] _134_\[8\] _06178_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__mux2_1
XFILLER_113_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11246_ _149_\[9\] _132_\[9\] VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__nand2_1
XFILLER_106_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11177_ _05227_ _05260_ _05261_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__a21o_1
XFILLER_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10128_ _01238_ _04032_ _04258_ _04500_ _01232_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__o311a_1
XFILLER_94_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10059_ _01244_ _03927_ _03929_ _04156_ _01238_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__a221o_1
XFILLER_94_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13818_ clknet_leaf_75_clk _01037_ VGND VGND VPWR VPWR _128_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13749_ clknet_leaf_75_clk _00968_ VGND VGND VPWR VPWR _132_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07270_ _182_\[5\] _01620_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__nand2_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09911_ _185_\[15\] _04150_ _04175_ _04293_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_7_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_113_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09842_ _185_\[12\] _04150_ _04175_ _04227_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__o211a_1
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _01230_ _03872_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__or2_1
XFILLER_86_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06985_ _243_\[25\] _01583_ _01557_ _01587_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__a211o_1
X_08724_ _03148_ _03149_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__nor2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08655_ _228_\[7\] _231_\[7\] _02790_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__a21oi_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07606_ _185_\[16\] _234_\[16\] VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__nand2_1
X_08586_ _228_\[5\] _231_\[5\] VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__nor2_1
XFILLER_42_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07537_ _01355_ _02080_ _02086_ _01884_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__a211o_1
XFILLER_35_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07468_ _01982_ _02005_ _02018_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__nand3_1
XFILLER_10_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07399_ _185_\[9\] _234_\[9\] VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__or2_1
XFILLER_6_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09207_ _02392_ _03617_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__or2_1
XFILLER_136_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09138_ _02327_ _03549_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__or2_1
XFILLER_135_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11100_ _158_\[1\] _158_\[0\] _05194_ _05196_ _158_\[2\] VGND VGND VPWR VPWR _05204_
+ sky130_fd_sc_hd__o311a_1
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09069_ _02842_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__xnor2_2
X_12080_ _140_\[2\] _142_\[2\] _06005_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__mux2_1
XFILLER_89_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11031_ _05159_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12982_ clknet_leaf_23_clk _00201_ VGND VGND VPWR VPWR _243_\[22\] sky130_fd_sc_hd__dfxtp_2
XFILLER_45_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11933_ _152_\[19\] _05933_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__nand2_1
XFILLER_91_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11864_ net4 _05776_ _05870_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__a22o_1
X_13603_ clknet_leaf_52_clk _00822_ VGND VGND VPWR VPWR _140_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10815_ _170_\[9\] _05002_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__or2_1
X_11795_ _01358_ _05808_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__and2_1
XFILLER_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13534_ clknet_leaf_66_clk _00753_ VGND VGND VPWR VPWR _152_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10746_ _170_\[21\] _173_\[21\] _04936_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__mux2_1
XFILLER_127_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13465_ clknet_leaf_123_clk _00684_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dfxtp_2
X_10677_ _01418_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__buf_2
X_12416_ _06242_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13396_ clknet_leaf_124_clk _00615_ VGND VGND VPWR VPWR _167_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12347_ _06206_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12278_ _136_\[0\] _134_\[0\] _06167_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__mux2_1
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11229_ _149_\[7\] _132_\[7\] VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__or2_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06770_ _179_\[1\] _01268_ _01251_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__or3_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08440_ _02842_ _02874_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__xnor2_2
XFILLER_90_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08371_ _02820_ _02791_ _02760_ _02821_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__o211a_1
X_07322_ _01802_ _01818_ _01850_ _01816_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__a211o_1
X_07253_ _01811_ _01812_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__or2_1
X_07184_ _01711_ _01739_ _01745_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__o21a_1
XFILLER_145_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09825_ _01242_ _03883_ _03984_ _04055_ _03876_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__a311o_1
XFILLER_86_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ _04114_ _04117_ _04143_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__o21a_1
XFILLER_104_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06968_ _243_\[20\] _01548_ _01545_ _01575_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__o211a_1
X_09687_ _03933_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__clkbuf_4
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08707_ _03132_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__inv_2
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ _01427_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__clkbuf_4
X_08638_ _170_\[6\] _02787_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__and2_1
XFILLER_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _02380_ _02977_ _02998_ _02999_ _01406_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__a221o_1
X_10600_ _173_\[8\] _176_\[8\] _01226_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__mux2_1
XFILLER_80_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11580_ _149_\[16\] _05615_ _05533_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__mux2_1
XFILLER_80_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10531_ _176_\[19\] _179_\[19\] _04790_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__mux2_1
X_13250_ clknet_leaf_8_clk _00469_ VGND VGND VPWR VPWR _182_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12201_ _06129_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__clkbuf_1
X_10462_ _04712_ _04764_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__or2_1
XFILLER_6_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10393_ _179_\[11\] _04684_ _04705_ _04715_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__o211a_1
X_13181_ clknet_leaf_102_clk _00400_ VGND VGND VPWR VPWR _225_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12132_ _06093_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12063_ _06038_ _06052_ _06042_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__a21o_1
XFILLER_89_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11014_ _04855_ _05148_ _05149_ _05122_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__a211o_1
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12965_ clknet_leaf_19_clk _00184_ VGND VGND VPWR VPWR _243_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11916_ _142_\[17\] _05918_ _05893_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__mux2_1
XFILLER_18_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12896_ clknet_leaf_72_clk _00120_ VGND VGND VPWR VPWR _116_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11847_ _140_\[21\] _05855_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__xnor2_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11778_ _152_\[5\] _05791_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__nor2_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13517_ clknet_leaf_80_clk _00736_ VGND VGND VPWR VPWR _152_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10729_ _170_\[16\] _04942_ _04922_ _04950_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__o211a_1
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13448_ clknet_leaf_2_clk _00667_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_2
XFILLER_126_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13379_ clknet_leaf_126_clk _00598_ VGND VGND VPWR VPWR _170_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07940_ _01354_ _02476_ _01412_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__o21ai_2
XFILLER_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07871_ _182_\[22\] _01678_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__or2_1
X_09610_ _01277_ _01279_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__and2b_1
X_06822_ _179_\[13\] _01300_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__or2_1
XFILLER_96_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09541_ _195_\[3\] _03874_ _195_\[0\] VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__or3b_2
XFILLER_95_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06753_ _179_\[0\] _01299_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__or2_1
XFILLER_55_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09472_ _03867_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__clkbuf_4
XFILLER_91_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06684_ _118_\[7\] _116_\[7\] _01370_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__mux2_1
XFILLER_70_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08423_ _225_\[28\] VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__buf_4
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08354_ _02749_ _02808_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__or2_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07305_ _01859_ _01862_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__xnor2_2
XFILLER_32_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08285_ _228_\[27\] _02733_ _02723_ _02756_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__o211a_1
XFILLER_20_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07236_ _01795_ _01796_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__xor2_1
XFILLER_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07167_ _01728_ _01729_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__nor2_1
XFILLER_145_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07098_ _01670_ _01673_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__or2_1
XFILLER_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09808_ _04153_ _04176_ _04193_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__o21bai_2
XFILLER_115_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09739_ _04120_ _04125_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__nor2_1
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12750_ _06417_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12681_ _06381_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11701_ _05722_ _05723_ _116_\[29\] VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11632_ _118_\[8\] _05661_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__xnor2_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13302_ clknet_leaf_8_clk _00521_ VGND VGND VPWR VPWR _176_\[16\] sky130_fd_sc_hd__dfxtp_1
X_11563_ _118_\[22\] _118_\[1\] VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11494_ _05522_ _05535_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__or2_1
X_10514_ _179_\[14\] _04799_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__or2_1
XFILLER_10_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13233_ clknet_leaf_25_clk _00452_ VGND VGND VPWR VPWR _182_\[11\] sky130_fd_sc_hd__dfxtp_1
X_10445_ _176_\[25\] _04725_ _04753_ _04728_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__a211o_1
XFILLER_109_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13164_ clknet_leaf_109_clk _00383_ VGND VGND VPWR VPWR _225_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12115_ _06084_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__clkbuf_1
X_10376_ _04692_ _04703_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__or2_1
X_13095_ clknet_leaf_106_clk _00314_ VGND VGND VPWR VPWR _231_\[7\] sky130_fd_sc_hd__dfxtp_1
X_12046_ _06037_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12948_ clknet_leaf_30_clk _00167_ VGND VGND VPWR VPWR _246_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _06484_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08070_ _02593_ _02601_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07021_ _01612_ _01565_ _01609_ _01613_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__o211a_1
XFILLER_115_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08972_ _02161_ _03348_ _03347_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__a21boi_2
X_07923_ _243_\[26\] _240_\[26\] _01690_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__mux2_4
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07854_ _02391_ _02392_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06805_ _246_\[8\] _01407_ _01436_ _01456_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__a211o_1
XFILLER_84_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07785_ _01698_ _02325_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__xnor2_2
XFILLER_45_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09524_ _246_\[1\] _01313_ _03913_ _243_\[1\] _01429_ VGND VGND VPWR VPWR _03921_
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06736_ _118_\[31\] _116_\[31\] _01394_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__mux2_1
XFILLER_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06667_ _01363_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09455_ _01923_ _03857_ _03858_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__or3_1
XFILLER_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08406_ _225_\[24\] VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__buf_4
X_06598_ _01300_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__clkbuf_2
X_09386_ _02549_ _03790_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__or2_1
XFILLER_137_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08337_ _02749_ _02795_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__or2_1
X_08268_ _231_\[22\] _02730_ _02712_ _02744_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__a211o_1
X_07219_ _01650_ _01632_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__xnor2_1
X_10230_ _01285_ _04107_ _04385_ _01239_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__o211a_1
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08199_ _01480_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10161_ _04532_ _04505_ _04506_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__a21o_1
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10092_ _04465_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__nor2_1
XFILLER_86_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13920_ clknet_leaf_70_clk _01139_ VGND VGND VPWR VPWR _120_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13851_ clknet_leaf_72_clk _01070_ VGND VGND VPWR VPWR _126_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12802_ _06444_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__clkbuf_1
X_13782_ clknet_leaf_94_clk _01001_ VGND VGND VPWR VPWR _130_\[22\] sky130_fd_sc_hd__dfxtp_1
X_10994_ _05079_ _05137_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__or2_1
X_12733_ _06408_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__clkbuf_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12664_ _06372_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__clkbuf_1
X_11615_ _116_\[20\] _05645_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__or2_1
X_12595_ _06336_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__clkbuf_1
X_11546_ _116_\[13\] _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__nor2_1
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13216_ clknet_leaf_37_clk _00435_ VGND VGND VPWR VPWR _185_\[26\] sky130_fd_sc_hd__dfxtp_4
X_11477_ _05501_ _05520_ _05522_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__o21ai_1
XFILLER_136_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10428_ _179_\[21\] _182_\[21\] _04693_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__mux2_1
XFILLER_124_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10359_ _04686_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__clkbuf_8
X_13147_ clknet_leaf_120_clk _00366_ VGND VGND VPWR VPWR _228_\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13078_ clknet_leaf_101_clk _00297_ VGND VGND VPWR VPWR _234_\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _06020_ _06021_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__or2_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07570_ _185_\[15\] _234_\[15\] VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__or2_1
XFILLER_53_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06521_ _195_\[5\] VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__buf_2
XFILLER_34_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09240_ _02431_ _03649_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09171_ _03581_ _03582_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__xor2_1
X_08122_ _234_\[12\] _02564_ _02629_ _02640_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__a211o_1
XFILLER_119_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08053_ _02584_ _02585_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__nor2_1
X_07004_ _243_\[31\] _01548_ _01598_ _01600_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__o211a_1
XFILLER_134_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08955_ _03273_ _03304_ _03336_ _03270_ _03303_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__o2111a_1
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07906_ _182_\[24\] _01684_ _02414_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__a21oi_2
XFILLER_57_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08886_ _02404_ _03306_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__nand2_1
XFILLER_84_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07837_ _02375_ _02376_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__nand2_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07768_ _02308_ _02309_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__or2_1
X_09507_ _01240_ _01283_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__or2_1
X_06719_ _01366_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__buf_4
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07699_ _185_\[19\] _234_\[19\] VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__or2_1
XFILLER_80_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09438_ _02380_ _03836_ _03842_ _01439_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__o211a_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09369_ _03765_ _03766_ _03775_ _01495_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__a211o_1
XFILLER_12_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11400_ _05452_ _05455_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__xnor2_1
X_12380_ _132_\[16\] _134_\[16\] _06219_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__mux2_1
XANTENNA_81 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11331_ _149_\[20\] _132_\[20\] VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__nand2_2
XANTENNA_70 _03568_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11262_ _149_\[11\] _132_\[11\] VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__nor2_1
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11193_ _149_\[2\] _132_\[2\] VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__nand2_1
X_10213_ _142_\[29\] _04581_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__and2_1
XFILLER_121_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13001_ clknet_leaf_20_clk _00220_ VGND VGND VPWR VPWR _240_\[9\] sky130_fd_sc_hd__dfxtp_1
X_10144_ _04513_ _04514_ _142_\[26\] VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_clk clknet_1_0_0_clk VGND VGND VPWR VPWR clknet_2_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_10075_ _04398_ _04404_ _04450_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__a21oi_2
XFILLER_102_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13903_ clknet_leaf_97_clk _01122_ VGND VGND VPWR VPWR _122_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13834_ clknet_leaf_93_clk _01053_ VGND VGND VPWR VPWR _126_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13765_ clknet_leaf_62_clk _00984_ VGND VGND VPWR VPWR _130_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10977_ net52 _05110_ _05126_ _05122_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__a211o_1
XFILLER_15_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13696_ clknet_leaf_59_clk _00915_ VGND VGND VPWR VPWR _134_\[0\] sky130_fd_sc_hd__dfxtp_1
X_12716_ _06399_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__clkbuf_1
X_12647_ _06363_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12578_ _06327_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__clkbuf_1
X_11529_ _05567_ _05569_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__nand2_1
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08740_ _03140_ _03142_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__and2b_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08671_ _03070_ _03085_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__nand2_1
XFILLER_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07622_ _182_\[16\] _01657_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__and2_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07553_ _02050_ _02076_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__or2_1
X_07484_ _02032_ _02034_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__nand2_1
X_06504_ _01216_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__buf_4
XFILLER_139_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09223_ _03630_ _03633_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__nand2_1
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09154_ _03499_ _03504_ _03534_ _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__a31o_1
X_08105_ _234_\[7\] _02448_ _02419_ _02628_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__o211a_1
X_09085_ _03428_ _03459_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__nand2_1
XFILLER_135_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08036_ _02557_ _02568_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__nor2_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09987_ _01292_ _04076_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__nor2_1
XFILLER_89_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08938_ _03354_ _03356_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08869_ _03288_ _03289_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__or2_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10900_ net47 _05048_ _05072_ _05067_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__o211a_1
XFILLER_29_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11880_ _152_\[14\] _05885_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__nand2_1
XFILLER_84_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10831_ _170_\[14\] _05002_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__or2_1
X_13550_ clknet_leaf_86_clk _00769_ VGND VGND VPWR VPWR _149_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10762_ _173_\[26\] _04953_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__or2_1
X_13481_ clknet_leaf_32_clk _00700_ _00114_ VGND VGND VPWR VPWR _190_\[3\] sky130_fd_sc_hd__dfrtp_1
X_12501_ _130_\[10\] _128_\[10\] _06280_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__mux2_1
XFILLER_40_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12432_ _132_\[9\] _130_\[9\] _06247_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__mux2_1
XFILLER_40_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10693_ _04671_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__clkbuf_4
X_12363_ _132_\[8\] _134_\[8\] _06208_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__mux2_1
XFILLER_138_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12294_ _01393_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__buf_4
XFILLER_107_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11314_ _05380_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__clkbuf_1
X_11245_ _149_\[9\] _132_\[9\] VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__nor2_1
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11176_ net24 _05190_ _05192_ _158_\[21\] VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__a22o_1
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10127_ _03979_ _04479_ _01238_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__o21ai_1
X_10058_ _04432_ _04433_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__or2_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13817_ clknet_leaf_71_clk _01036_ VGND VGND VPWR VPWR _128_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13748_ clknet_leaf_77_clk _00967_ VGND VGND VPWR VPWR _132_\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_44_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13679_ clknet_leaf_78_clk _00898_ VGND VGND VPWR VPWR _136_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09910_ _04289_ _04291_ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__o21ai_1
X_09841_ _04225_ _04226_ _03946_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__a21o_1
XFILLER_113_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _04075_ _03897_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__nor2_1
X_06984_ _240_\[25\] _01565_ _01558_ _01586_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__o211a_1
XFILLER_58_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _228_\[9\] _231_\[9\] _02797_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__a21oi_2
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08654_ _228_\[7\] _231_\[7\] VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__nor2_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _03012_ _03014_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__xnor2_2
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07605_ _185_\[16\] _234_\[16\] VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__or2_1
X_07536_ _01778_ _02085_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__nor2_1
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07467_ _01982_ _02005_ _02018_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__a21oi_1
X_09206_ _03615_ _03616_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__and2_1
XFILLER_22_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07398_ _01671_ _01951_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__xnor2_1
X_09137_ _02327_ _03549_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__nand2_1
XFILLER_136_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09068_ _02801_ _02772_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08019_ _02511_ _02538_ _02550_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__nor3_1
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11030_ _01710_ _05158_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__or2_1
XFILLER_134_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12981_ clknet_leaf_23_clk _00200_ VGND VGND VPWR VPWR _243_\[21\] sky130_fd_sc_hd__dfxtp_2
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11932_ _140_\[29\] _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__xnor2_2
XFILLER_17_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11863_ _05864_ _05869_ _05785_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__o21a_1
XFILLER_72_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13602_ clknet_leaf_52_clk _00821_ VGND VGND VPWR VPWR _140_\[2\] sky130_fd_sc_hd__dfxtp_2
X_10814_ _164_\[8\] _04986_ _05011_ _05001_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__a211o_1
XFILLER_32_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11794_ _05793_ _05806_ _05801_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__or3_1
XFILLER_13_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13533_ clknet_leaf_67_clk _00752_ VGND VGND VPWR VPWR _152_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10745_ _167_\[20\] _04925_ _04962_ _04939_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__o211a_1
XFILLER_43_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10676_ _170_\[1\] _04833_ _04806_ _04912_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__o211a_1
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13464_ clknet_leaf_123_clk _00683_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dfxtp_2
X_12415_ _132_\[1\] _130_\[1\] _06201_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__mux2_1
X_13395_ clknet_leaf_124_clk _00614_ VGND VGND VPWR VPWR _167_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12346_ _132_\[0\] _134_\[0\] _06090_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__mux2_1
XFILLER_5_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12277_ _06169_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11228_ _05305_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11159_ _158_\[16\] _01262_ _158_\[17\] VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08370_ net43 _02798_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__or2_1
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07321_ _01877_ _01878_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__nor2_1
XFILLER_32_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07252_ _01782_ _01804_ _01810_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__and3_1
XFILLER_136_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07183_ _182_\[1\] _01604_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__nand2_1
XFILLER_145_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_815 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09824_ _03910_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09755_ _04114_ _04117_ _04143_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__or3_1
XFILLER_74_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06967_ _01568_ _01574_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__or2_1
XFILLER_73_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09686_ _03923_ _04076_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__nor2_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06898_ _243_\[0\] _01496_ _01509_ _01525_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__a211o_1
X_08706_ _03130_ _03131_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__xnor2_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08637_ _03063_ _03064_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__nor2_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _02964_ _02997_ _02996_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07519_ _02064_ _02067_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__nand2_1
X_08499_ _170_\[0\] _02768_ _02906_ _02931_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__a31oi_4
X_10530_ _173_\[18\] _04774_ _04813_ _04777_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__a211o_1
XFILLER_109_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10461_ _179_\[31\] _182_\[31\] _04743_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__mux2_1
XFILLER_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12200_ _140_\[27\] _138_\[27\] _06123_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__mux2_1
XFILLER_136_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10392_ _182_\[11\] _04696_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__or2_1
X_13180_ clknet_leaf_102_clk _00399_ VGND VGND VPWR VPWR _225_\[28\] sky130_fd_sc_hd__dfxtp_1
X_12131_ _140_\[26\] _142_\[26\] _06090_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__mux2_1
XFILLER_89_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12062_ _06041_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__inv_2
XFILLER_104_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11013_ _03060_ _04631_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__nor2_1
XFILLER_89_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12964_ clknet_leaf_20_clk _00183_ VGND VGND VPWR VPWR _243_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11915_ net9 _05917_ _05852_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__mux2_1
X_12895_ clknet_leaf_72_clk _00119_ VGND VGND VPWR VPWR _116_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11846_ _140_\[28\] _140_\[30\] VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__xnor2_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11777_ _152_\[5\] _05791_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__nand2_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13516_ clknet_leaf_78_clk _00735_ VGND VGND VPWR VPWR _152_\[12\] sky130_fd_sc_hd__dfxtp_1
X_10728_ _173_\[16\] _04917_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__or2_1
XFILLER_41_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10659_ _02483_ _04691_ _04901_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__o21a_1
X_13447_ clknet_leaf_12_clk _00666_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dfxtp_4
XFILLER_127_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13378_ clknet_leaf_127_clk _00597_ VGND VGND VPWR VPWR _170_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12329_ _06196_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07870_ _02351_ _02408_ _02297_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__o21a_1
XFILLER_110_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06821_ _246_\[12\] _01422_ _01425_ _01468_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__o211a_1
XFILLER_56_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09540_ _01240_ _03935_ _03936_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__or3_1
XFILLER_110_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06752_ _01411_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__clkbuf_4
XFILLER_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09471_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__buf_2
XFILLER_83_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06683_ _01373_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08422_ _02711_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08353_ net39 _02807_ _02750_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__mux2_1
X_07304_ _01822_ _01823_ _01860_ _01829_ _01861_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__o311a_1
X_08284_ _164_\[27\] _02736_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__or2_1
X_07235_ _01736_ _01765_ _01764_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__a21bo_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07166_ _185_\[1\] _234_\[1\] VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__nor2_1
XFILLER_132_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07097_ _173_\[20\] _01671_ _01672_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__mux2_1
XFILLER_121_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09807_ _04153_ _04176_ _04193_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__or3b_1
XFILLER_101_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07999_ _02532_ _02533_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__or2b_1
X_09738_ _185_\[8\] _03869_ _03919_ _04127_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__o211a_1
XFILLER_115_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09669_ _01292_ _04057_ _04059_ _04060_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__o211a_1
XFILLER_82_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12680_ _126_\[31\] _124_\[31\] _06379_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__mux2_1
X_11700_ _118_\[4\] _118_\[15\] VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__nand2_1
XFILLER_70_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _118_\[25\] _118_\[29\] VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__xnor2_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11562_ _05599_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10513_ _173_\[13\] _04774_ _04801_ _04777_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__a211o_1
X_13301_ clknet_leaf_25_clk _00520_ VGND VGND VPWR VPWR _176_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11493_ _05517_ _05528_ _05529_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__o21a_1
XFILLER_6_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13232_ clknet_leaf_27_clk _00451_ VGND VGND VPWR VPWR _182_\[10\] sky130_fd_sc_hd__dfxtp_1
X_10444_ _179_\[25\] _04721_ _04751_ _04752_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__o211a_1
XFILLER_108_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10375_ _179_\[6\] _182_\[6\] _04693_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__mux2_1
X_13163_ clknet_leaf_106_clk _00382_ VGND VGND VPWR VPWR _225_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12114_ _140_\[18\] _142_\[18\] _06079_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__mux2_1
XFILLER_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13094_ clknet_leaf_111_clk _00313_ VGND VGND VPWR VPWR _231_\[6\] sky130_fd_sc_hd__dfxtp_1
X_12045_ _142_\[28\] _06036_ _06005_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__mux2_1
XFILLER_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12947_ clknet_leaf_30_clk _00166_ VGND VGND VPWR VPWR _246_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _118_\[30\] _120_\[30\] _01361_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__mux2_1
XFILLER_61_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11829_ _05823_ _05830_ _05838_ _01274_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__a31o_1
XFILLER_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07020_ _173_\[3\] _01580_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__or2_1
XFILLER_142_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08971_ _02192_ _03388_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07922_ _02457_ _02458_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__or2_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07853_ _243_\[24\] _240_\[24\] _01684_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__mux2_4
X_06804_ _243_\[8\] _01438_ _01439_ _01455_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__o211a_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07784_ _01654_ _01604_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09523_ _142_\[0\] _03915_ _03916_ _03912_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__o2bb2ai_1
X_06735_ _01401_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06666_ _116_\[0\] _118_\[0\] _01362_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__mux2_1
X_09454_ _03832_ _03844_ _03856_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08405_ _228_\[23\] _02845_ _02834_ _02848_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__o211a_1
X_09385_ _02549_ _03790_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__nand2_1
X_06597_ _01299_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__clkbuf_2
XFILLER_101_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08336_ net66 _02794_ _02750_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__mux2_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08267_ _228_\[22\] _02733_ _02723_ _02743_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__o211a_1
XFILLER_20_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07218_ _01755_ _01756_ _01757_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__nand3_1
X_08198_ _231_\[2\] _02659_ _02636_ _02694_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__o211a_1
X_07149_ _01638_ _01623_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10160_ _04486_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__inv_2
XFILLER_105_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10091_ _04432_ _04444_ _04464_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__o21a_1
XFILLER_87_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13850_ clknet_leaf_89_clk _01069_ VGND VGND VPWR VPWR _126_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12801_ _122_\[25\] _120_\[25\] _06434_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__mux2_1
X_13781_ clknet_leaf_93_clk _01000_ VGND VGND VPWR VPWR _130_\[21\] sky130_fd_sc_hd__dfxtp_1
X_10993_ _164_\[30\] _167_\[30\] _01214_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__mux2_1
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12732_ _124_\[24\] _122_\[24\] _06401_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__mux2_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12663_ _126_\[23\] _124_\[23\] _06368_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__mux2_1
XFILLER_128_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11614_ _116_\[20\] _05645_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__nand2_1
X_12594_ _128_\[22\] _126_\[22\] _06335_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__mux2_1
XFILLER_11_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11545_ _118_\[20\] _05583_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__xnor2_1
X_11476_ _116_\[5\] _05510_ _05521_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__o21ai_1
XFILLER_7_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13215_ clknet_leaf_37_clk _00434_ VGND VGND VPWR VPWR _185_\[25\] sky130_fd_sc_hd__dfxtp_4
XFILLER_109_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10427_ _176_\[20\] _04735_ _04739_ _04740_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__o211a_1
XFILLER_7_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10358_ _176_\[1\] _04683_ _04690_ _01419_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__a211o_1
X_13146_ clknet_leaf_120_clk _00365_ VGND VGND VPWR VPWR _228_\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10289_ _01423_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__clkbuf_8
X_13077_ clknet_leaf_100_clk _00296_ VGND VGND VPWR VPWR _234_\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12028_ _06018_ _06019_ _152_\[27\] VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13979_ clknet_leaf_90_clk _01198_ VGND VGND VPWR VPWR _118_\[27\] sky130_fd_sc_hd__dfxtp_2
XFILLER_53_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06520_ _01229_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09170_ _03550_ _03551_ _03553_ _03554_ _02337_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__a32o_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08121_ _231_\[12\] _02611_ _01695_ _02639_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_122_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_122_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_107_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08052_ _02546_ _02571_ _02583_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__nor3_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07003_ _01568_ _01599_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__or2_1
XFILLER_1_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08954_ _170_\[15\] _02817_ _02814_ _170_\[14\] VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__o211a_1
X_07905_ _02441_ _02442_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__nand2_1
XFILLER_96_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08885_ _03303_ _03305_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__xor2_2
XFILLER_84_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07836_ _02341_ _02345_ _02339_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__a21bo_1
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07767_ _02264_ _02265_ _02307_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__and3_1
X_09506_ _03901_ _03903_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__nand2_1
X_06718_ _01391_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07698_ _02241_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__inv_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06649_ _01295_ _01324_ _01349_ _01272_ _01307_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__o2111a_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09437_ _02404_ _03841_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__nand2_1
XFILLER_9_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09368_ _01437_ _03774_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__and2_1
XFILLER_12_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08319_ net62 _02781_ _02750_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_113_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_113_clk sky130_fd_sc_hd__clkbuf_16
X_09299_ _03685_ _03687_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__and2b_1
XANTENNA_71 _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ _149_\[20\] _132_\[20\] VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__or2_1
XANTENNA_60 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11261_ _05279_ _05331_ _05333_ _05334_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__a31o_1
XFILLER_125_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11192_ _149_\[2\] _132_\[2\] VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__nor2_1
X_10212_ _246_\[29\] _01316_ _04409_ _243_\[29\] _01513_ VGND VGND VPWR VPWR _04581_
+ sky130_fd_sc_hd__o221a_1
X_13000_ clknet_leaf_19_clk _00219_ VGND VGND VPWR VPWR _240_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10143_ _142_\[26\] _04513_ _04514_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__and3_1
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10074_ _04395_ _04425_ _04426_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__or3b_1
XFILLER_48_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13902_ clknet_leaf_98_clk _01121_ VGND VGND VPWR VPWR _122_\[14\] sky130_fd_sc_hd__dfxtp_1
X_13833_ clknet_leaf_62_clk _01052_ VGND VGND VPWR VPWR _126_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13764_ clknet_leaf_62_clk _00983_ VGND VGND VPWR VPWR _130_\[4\] sky130_fd_sc_hd__dfxtp_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10976_ _164_\[24\] _05107_ _05094_ _05125_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__o211a_1
X_13695_ clknet_leaf_58_clk _00914_ VGND VGND VPWR VPWR _136_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12715_ _124_\[16\] _122_\[16\] _06390_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__mux2_1
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12646_ _126_\[15\] _124_\[15\] _06357_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_104_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_104_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_117_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12577_ _128_\[14\] _126_\[14\] _06324_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__mux2_1
XFILLER_144_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11528_ _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__inv_2
X_11459_ _05501_ _05506_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__xor2_1
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ clknet_leaf_117_clk _00348_ VGND VGND VPWR VPWR _228_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_787 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08670_ _03050_ _03086_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__nand2_1
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07621_ _182_\[16\] _01657_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__nor2_1
X_07552_ _02098_ _02100_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06503_ _01212_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__clkbuf_4
X_07483_ _01962_ _01992_ _02031_ _02033_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__a31oi_2
XFILLER_34_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09222_ _03503_ _03631_ _03629_ _03632_ _03368_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__o32a_1
X_09153_ _03565_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__inv_2
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08104_ _02625_ _02627_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__or2_1
X_09084_ _03497_ _03498_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__and2_1
X_08035_ _02531_ _02532_ _02533_ _02558_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__o211a_1
XFILLER_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09986_ _04010_ _03952_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__and2b_1
XFILLER_107_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08937_ _228_\[16\] _231_\[16\] _03355_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__o21a_1
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08868_ _03285_ _03287_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__and2_1
XFILLER_57_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07819_ _02357_ _02358_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__xnor2_4
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08799_ _185_\[12\] _03221_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10830_ _01225_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__clkbuf_4
X_10761_ _167_\[25\] _04925_ _04973_ _04939_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__o211a_1
XFILLER_13_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12500_ _06286_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__clkbuf_1
X_13480_ clknet_leaf_28_clk _00699_ _00113_ VGND VGND VPWR VPWR _190_\[2\] sky130_fd_sc_hd__dfrtp_1
X_10692_ _167_\[5\] _04836_ _04924_ _04914_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__a211o_1
XFILLER_40_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12431_ _06250_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12362_ _06214_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12293_ _06177_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__clkbuf_1
X_11313_ _152_\[17\] _05379_ _05318_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__mux2_1
X_11244_ _05319_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11175_ _01266_ _05259_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__nand2_1
XFILLER_68_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10126_ _04438_ _04498_ _01238_ _04365_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_79_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10057_ _142_\[22\] _04431_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__nor2_1
XFILLER_94_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13816_ clknet_leaf_68_clk _01035_ VGND VGND VPWR VPWR _128_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13747_ clknet_leaf_74_clk _00966_ VGND VGND VPWR VPWR _132_\[19\] sky130_fd_sc_hd__dfxtp_1
X_10959_ _05079_ _05113_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__or2_1
XFILLER_16_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13678_ clknet_leaf_47_clk _00897_ VGND VGND VPWR VPWR _136_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12629_ _126_\[7\] _124_\[7\] _06346_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__mux2_1
XFILLER_129_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09840_ _04205_ _04224_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__nand2_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _04156_ _03925_ _04157_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__a211o_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06983_ _176_\[25\] _01580_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__or2_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _228_\[9\] _231_\[9\] VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__nor2_1
XFILLER_54_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08653_ _03078_ _03080_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__xnor2_2
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08584_ _01814_ _02986_ _03013_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__a21oi_2
X_07604_ _02150_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__inv_2
XFILLER_42_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07535_ _02083_ _02084_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__xnor2_2
X_07466_ _02016_ _02017_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__xor2_1
XFILLER_50_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09205_ _03608_ _03610_ _03614_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__nand3_1
X_07397_ _01654_ _01608_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09136_ _185_\[22\] _03548_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__xnor2_1
X_09067_ _02252_ _03449_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__nand2_1
X_08018_ _02551_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__inv_2
XFILLER_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09969_ _04327_ _04328_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nor2_1
XFILLER_103_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12980_ clknet_leaf_23_clk _00199_ VGND VGND VPWR VPWR _243_\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11931_ _140_\[4\] _140_\[6\] VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__xnor2_2
XFILLER_45_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11862_ _05864_ _05869_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__nand2_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13601_ clknet_leaf_53_clk _00820_ VGND VGND VPWR VPWR _140_\[1\] sky130_fd_sc_hd__dfxtp_2
X_10813_ _167_\[8\] _04980_ _05009_ _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__o211a_1
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11793_ _05793_ _05801_ _05806_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__o21ai_1
X_13532_ clknet_leaf_67_clk _00751_ VGND VGND VPWR VPWR _152_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10744_ _04888_ _04961_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__or2_1
X_10675_ _173_\[1\] _04799_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__or2_1
X_13463_ clknet_leaf_1_clk _00682_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfxtp_4
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12414_ _06241_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__clkbuf_1
X_13394_ clknet_leaf_124_clk _00613_ VGND VGND VPWR VPWR _167_\[12\] sky130_fd_sc_hd__dfxtp_1
X_12345_ _06205_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12276_ _138_\[31\] _136_\[31\] _06167_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__mux2_1
XFILLER_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11227_ _152_\[6\] _05304_ _01362_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__mux2_1
X_11158_ _05227_ _05246_ _05247_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__a21o_1
X_10109_ _04477_ _04478_ _04481_ _04474_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__o31a_1
XFILLER_110_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11089_ net35 _01325_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__or2_1
XFILLER_83_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07320_ _01844_ _01865_ _01876_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__nor3_1
X_07251_ _01782_ _01804_ _01810_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__a21oi_1
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07182_ _01744_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09823_ _04207_ _04208_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__nor2_1
XFILLER_99_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09754_ _04131_ _04142_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__xor2_1
X_06966_ _176_\[20\] _240_\[20\] _01569_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__mux2_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09685_ _04002_ _01278_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__or2_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06897_ _240_\[0\] _01474_ _01510_ _01524_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__o211a_1
XFILLER_67_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08705_ _03122_ _03121_ _03123_ _03120_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__a31oi_2
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_93_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_16
X_08636_ _170_\[7\] _02790_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__and2_1
XFILLER_27_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08567_ _02964_ _02996_ _02997_ _01523_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__o31a_1
X_07518_ _02064_ _02067_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__or2_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08498_ _170_\[1\] _02772_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__and2_1
X_07449_ _01404_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__clkbuf_4
X_10460_ _176_\[30\] _04735_ _04763_ _04740_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__o211a_1
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09119_ _03491_ _03513_ _03531_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__or3_1
XFILLER_129_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10391_ _176_\[10\] _04691_ _04714_ _04677_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__o211a_1
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12130_ _06092_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12061_ _06049_ _06050_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__nand2_1
XFILLER_89_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11012_ net64 _164_\[6\] _01215_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__mux2_1
XFILLER_2_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12963_ clknet_leaf_40_clk _00182_ VGND VGND VPWR VPWR _243_\[3\] sky130_fd_sc_hd__dfxtp_1
X_11914_ _05915_ _05916_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_84_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_18_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12894_ clknet_leaf_71_clk _00118_ VGND VGND VPWR VPWR _116_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11845_ _05854_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__clkbuf_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11776_ _140_\[22\] _05790_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__xnor2_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13515_ clknet_leaf_81_clk _00734_ VGND VGND VPWR VPWR _152_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10727_ _167_\[15\] _04945_ _04949_ _04914_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__a211o_1
X_13446_ clknet_leaf_123_clk _00665_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_2
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10658_ _176_\[27\] _04678_ _04633_ _173_\[27\] _04648_ VGND VGND VPWR VPWR _04901_
+ sky130_fd_sc_hd__o221a_1
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10589_ _04630_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__buf_4
X_13377_ clknet_leaf_127_clk _00596_ VGND VGND VPWR VPWR _170_\[27\] sky130_fd_sc_hd__dfxtp_2
XFILLER_115_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12328_ _136_\[24\] _134_\[24\] _06189_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__mux2_1
XFILLER_141_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12259_ _138_\[23\] _136_\[23\] _06156_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__mux2_1
XFILLER_5_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06820_ _01444_ _01467_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__nand2_1
XFILLER_95_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06751_ _01410_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__buf_6
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09470_ _03867_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_75_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_16
X_06682_ _118_\[6\] _116_\[6\] _01370_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__mux2_1
XFILLER_36_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08421_ _228_\[27\] _02838_ _02810_ _02860_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__a211o_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08352_ _225_\[12\] VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__clkbuf_4
X_07303_ _182_\[4\] _01616_ _01828_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__nand3_1
X_08283_ _231_\[26\] _02730_ _02753_ _02755_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__a211o_1
XFILLER_20_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07234_ _01793_ _01794_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__nand2_1
XFILLER_118_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07165_ _185_\[1\] _234_\[1\] VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__and2_1
XFILLER_145_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07096_ _01518_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__buf_4
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09806_ _04191_ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__or2_1
XFILLER_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07998_ _182_\[28\] _01698_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__nand2_1
X_09737_ _04125_ _04126_ _03868_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__o21ai_1
XFILLER_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06949_ _240_\[15\] _01526_ _01558_ _01561_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_66_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_16
X_09668_ _01230_ _01235_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__nor2_2
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09599_ _03992_ _03993_ _03946_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__a21o_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _03044_ _03047_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__xnor2_2
XFILLER_54_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11630_ _05659_ _05660_ _149_\[21\] _05262_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11561_ _149_\[14\] _05598_ _05533_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__mux2_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10512_ _176_\[13\] _04771_ _04751_ _04800_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__o211a_1
X_13300_ clknet_leaf_9_clk _00519_ VGND VGND VPWR VPWR _176_\[14\] sky130_fd_sc_hd__dfxtp_1
X_11492_ _05520_ _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__or2_1
XFILLER_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13231_ clknet_leaf_27_clk _00450_ VGND VGND VPWR VPWR _182_\[9\] sky130_fd_sc_hd__dfxtp_1
X_10443_ _182_\[25\] _04746_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__or2_1
XFILLER_40_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10374_ _176_\[5\] _04683_ _04702_ _01419_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__a211o_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13162_ clknet_leaf_106_clk _00381_ VGND VGND VPWR VPWR _225_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12113_ _06083_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13093_ clknet_leaf_111_clk _00312_ VGND VGND VPWR VPWR _231_\[5\] sky130_fd_sc_hd__dfxtp_1
X_12044_ net21 _06035_ _05785_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__mux2_1
XFILLER_77_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12946_ clknet_leaf_21_clk _00165_ VGND VGND VPWR VPWR _246_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _06483_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__clkbuf_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _05823_ _05830_ _05838_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__a21oi_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11759_ _05775_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13429_ clknet_leaf_123_clk _00648_ VGND VGND VPWR VPWR _164_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08970_ _03385_ _03387_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__xor2_1
XFILLER_130_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07921_ _02424_ _02425_ _02456_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__and3_1
XFILLER_96_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07852_ _02389_ _02390_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__or2_1
XFILLER_29_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06803_ _179_\[8\] _01299_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__or2_1
XFILLER_84_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 din[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_09522_ _02833_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_48_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_83_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07783_ _02323_ _02306_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__or2_1
X_06734_ _118_\[30\] _116_\[30\] _01394_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__mux2_1
XFILLER_71_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06665_ _01361_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__buf_4
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09453_ _03832_ _03844_ _03856_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__and3_1
XFILLER_37_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08404_ _02002_ _02847_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__or2_1
X_09384_ _03788_ _03789_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__and2_1
X_06596_ _01268_ _01251_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__or2_2
X_08335_ _225_\[8\] VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__buf_4
XFILLER_138_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08266_ _164_\[22\] _02736_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__or2_1
XFILLER_20_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07217_ _01353_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__clkbuf_4
X_08197_ _02686_ _02693_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__or2_1
XFILLER_106_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07148_ _182_\[0\] _237_\[0\] VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__or2_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07079_ _01657_ _01639_ _01609_ _01658_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__o211a_1
XFILLER_133_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10090_ _04432_ _04444_ _04464_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__nor3_1
XFILLER_114_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_74_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12800_ _06443_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13780_ clknet_leaf_93_clk _00999_ VGND VGND VPWR VPWR _130_\[20\] sky130_fd_sc_hd__dfxtp_1
X_10992_ net57 _05110_ _05136_ _05122_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__a211o_1
XFILLER_55_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12731_ _06407_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12662_ _06371_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__clkbuf_1
X_11613_ _118_\[6\] _05644_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__xnor2_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12593_ _06200_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__buf_4
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11544_ _118_\[16\] _118_\[31\] VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11475_ _116_\[4\] _05503_ _05510_ _116_\[5\] VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__a22o_1
XFILLER_137_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13214_ clknet_leaf_37_clk _00433_ VGND VGND VPWR VPWR _185_\[24\] sky130_fd_sc_hd__dfxtp_4
XFILLER_109_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10426_ _01424_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10357_ _179_\[1\] _04684_ _04686_ _04689_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__o211a_1
X_13145_ clknet_leaf_119_clk _00364_ VGND VGND VPWR VPWR _228_\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10288_ _179_\[7\] _04646_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__or2_1
XFILLER_78_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13076_ clknet_leaf_99_clk _00295_ VGND VGND VPWR VPWR _234_\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12027_ _152_\[27\] _06018_ _06019_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__and3_1
XFILLER_78_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13978_ clknet_leaf_91_clk _01197_ VGND VGND VPWR VPWR _118_\[26\] sky130_fd_sc_hd__dfxtp_2
XFILLER_46_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12929_ clknet_leaf_41_clk _00148_ VGND VGND VPWR VPWR _246_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08120_ _167_\[12\] _02616_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__or2_1
XFILLER_135_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08051_ _02546_ _02571_ _02583_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__o21a_1
XFILLER_134_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07002_ _176_\[31\] _240_\[31\] _01569_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__mux2_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08953_ _03370_ _03371_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__nand2_2
X_07904_ _182_\[25\] _01687_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__or2_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08884_ _03273_ _03304_ _03270_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__o21ai_2
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07835_ _02373_ _02374_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__and2b_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07766_ _02264_ _02265_ _02307_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__a21oi_1
X_09505_ _03902_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__clkbuf_4
X_06717_ _118_\[23\] _116_\[23\] _01381_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__mux2_1
XFILLER_80_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07697_ _01704_ _02240_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__xnor2_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ _03839_ _03840_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__xor2_2
XFILLER_25_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06648_ _01250_ _01207_ _01208_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__or3b_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06579_ _01233_ _01287_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09367_ _03770_ _03773_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__xnor2_1
XANTENNA_50 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08318_ _225_\[4\] VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__clkbuf_4
X_09298_ _02855_ _01426_ _03379_ _03706_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__o211a_1
XANTENNA_72 _04577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08249_ _164_\[17\] _02701_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__or2_1
XANTENNA_83 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11260_ _152_\[10\] _01368_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__and2_1
XFILLER_118_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10211_ _04574_ _04575_ _04577_ _04579_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__o2bb2a_1
X_11191_ _05264_ _05268_ _05272_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__o21a_1
XFILLER_106_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10142_ _246_\[26\] _01316_ _01301_ _179_\[26\] VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__o22a_1
XFILLER_121_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10073_ _04447_ _04448_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__and2_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13901_ clknet_leaf_97_clk _01120_ VGND VGND VPWR VPWR _122_\[13\] sky130_fd_sc_hd__dfxtp_1
X_13832_ clknet_leaf_62_clk _01051_ VGND VGND VPWR VPWR _126_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13763_ clknet_leaf_63_clk _00982_ VGND VGND VPWR VPWR _130_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10975_ _167_\[24\] _04867_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__or2_1
X_12714_ _06398_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__clkbuf_1
X_13694_ clknet_leaf_58_clk _00913_ VGND VGND VPWR VPWR _136_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12645_ _06362_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12576_ _06326_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__clkbuf_1
X_11527_ _116_\[11\] _05566_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__nor2_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11458_ _05504_ _05505_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__nand2_1
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11389_ _05434_ _05442_ _05445_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__o21ai_1
X_10409_ _01418_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__clkbuf_4
XFILLER_98_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13128_ clknet_leaf_111_clk _00347_ VGND VGND VPWR VPWR _228_\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13059_ clknet_leaf_15_clk _00278_ VGND VGND VPWR VPWR _234_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07620_ _02148_ _02165_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__or2_1
X_07551_ _02070_ _02072_ _02099_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__o21ba_1
X_06502_ _01215_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_6
X_07482_ _01986_ _01988_ _02020_ _02019_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__a31o_1
X_09221_ _03501_ _03631_ _03629_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__or3_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09152_ _03497_ _03532_ _03533_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__a21bo_1
X_08103_ _167_\[7\] _231_\[7\] _02626_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__mux2_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09083_ _03479_ _03480_ _03496_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__or3_1
XFILLER_135_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08034_ _02565_ _02566_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__nand2_1
XFILLER_143_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09985_ _03896_ _04132_ _04363_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__a21oi_1
XFILLER_103_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08936_ _228_\[16\] _231_\[16\] _02820_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__a21o_1
XFILLER_97_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08867_ _03285_ _03287_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__nor2_1
XFILLER_84_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07818_ _02350_ _02352_ _02349_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__a21oi_2
XFILLER_45_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08798_ _02852_ _03220_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__xnor2_2
X_07749_ _02290_ _02285_ _02287_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__and3_1
XFILLER_37_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10760_ _04971_ _04972_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__or2_1
XFILLER_52_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10691_ _170_\[5\] _04833_ _04922_ _04923_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__o211a_1
X_09419_ _02582_ _03823_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__xnor2_1
X_12430_ _132_\[8\] _130_\[8\] _06247_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__mux2_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12361_ _132_\[7\] _134_\[7\] _06208_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__mux2_1
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12292_ _136_\[7\] _134_\[7\] _06167_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__mux2_1
X_11312_ _05377_ _05378_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__xnor2_1
X_11243_ _152_\[8\] _05317_ _05318_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__mux2_1
XFILLER_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11174_ _158_\[21\] _01265_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__nand2_1
X_10125_ _03887_ _03925_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__nand2_1
XFILLER_121_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10056_ _142_\[22\] _04431_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__and2_1
XFILLER_102_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13815_ clknet_leaf_93_clk _01034_ VGND VGND VPWR VPWR _128_\[23\] sky130_fd_sc_hd__dfxtp_1
X_13746_ clknet_leaf_74_clk _00965_ VGND VGND VPWR VPWR _132_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10958_ _164_\[19\] _167_\[19\] _05064_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__mux2_1
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13677_ clknet_leaf_78_clk _00896_ VGND VGND VPWR VPWR _136_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12628_ _06353_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__clkbuf_1
X_10889_ _01213_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__buf_4
XFILLER_12_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12559_ _06317_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09770_ _03934_ _04005_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__nor2_1
XFILLER_98_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06982_ _243_\[24\] _01583_ _01557_ _01585_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__a211o_1
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08721_ _03144_ _03146_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__xnor2_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ _01875_ _03040_ _03079_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__a21oi_2
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07603_ _01694_ _02149_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08583_ _02983_ _02985_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__and2b_1
X_07534_ _182_\[12\] _01642_ _02056_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07465_ _243_\[11\] _240_\[11\] _01638_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__mux2_2
XFILLER_22_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09204_ _03608_ _03610_ _03614_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__a21o_1
X_07396_ _01938_ _01939_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__and2b_1
XFILLER_136_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09135_ _02849_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__xnor2_2
X_09066_ _03446_ _03448_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__or2b_1
XFILLER_135_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08017_ _02511_ _02538_ _02550_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__o21ai_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09968_ _04327_ _04328_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__nand2_1
XFILLER_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08919_ _01409_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__nand2_1
X_09899_ _03888_ _04006_ _04080_ _01243_ _01237_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__a221o_1
X_11930_ _05931_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11861_ _05867_ _05868_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__nand2_1
XFILLER_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11792_ _05804_ _05805_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__nand2_1
X_13600_ clknet_leaf_53_clk _00819_ VGND VGND VPWR VPWR _140_\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_60_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10812_ _170_\[8\] _05002_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__or2_1
XFILLER_13_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13531_ clknet_leaf_67_clk _00750_ VGND VGND VPWR VPWR _152_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10743_ _170_\[20\] _173_\[20\] _04936_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__mux2_1
XFILLER_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13462_ clknet_leaf_123_clk _00681_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfxtp_4
X_10674_ _167_\[0\] _04818_ _04911_ _04891_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__o211a_1
X_12413_ _132_\[0\] _130_\[0\] _06201_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__mux2_1
X_13393_ clknet_leaf_130_clk _00612_ VGND VGND VPWR VPWR _167_\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_138_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12344_ _136_\[31\] _134_\[31\] _06201_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__mux2_1
XFILLER_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12275_ _06168_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__clkbuf_1
X_11226_ _05301_ _05303_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__xor2_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11157_ net18 _05202_ _05193_ _158_\[16\] VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__a22o_1
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10108_ _04474_ _04477_ _04478_ _04481_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__nor4_1
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11088_ _01303_ _01318_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__nand2_4
XFILLER_76_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10039_ _01244_ _03928_ _03929_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__and3_1
XFILLER_48_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13729_ clknet_leaf_57_clk _00948_ VGND VGND VPWR VPWR _132_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07250_ _01806_ _01809_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__xor2_1
XFILLER_32_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07181_ _01710_ _01743_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__or2_1
XFILLER_117_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09822_ _142_\[12\] _04206_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__nor2_1
XFILLER_86_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09753_ _04134_ _04136_ _04141_ _01231_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__a22o_1
XFILLER_98_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06965_ _243_\[19\] _01548_ _01545_ _01573_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__o211a_1
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ _03128_ _03129_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__nand2_1
X_09684_ _04002_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__buf_2
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06896_ _176_\[0\] _01523_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__or2_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08635_ _170_\[7\] _02790_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__nor2_1
XFILLER_82_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _02967_ _02965_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__nor2_1
XFILLER_42_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07517_ _02065_ _02066_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__nand2_1
X_08497_ _02904_ _02928_ _01302_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__o21a_1
X_07448_ _01998_ _02000_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__xor2_2
XFILLER_109_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07379_ _01933_ _01934_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__nand2_1
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09118_ _03491_ _03513_ _03531_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__o21ai_1
XFILLER_108_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10390_ _04712_ _04713_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__or2_1
XFILLER_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09049_ _01409_ _03464_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__nand2_1
XFILLER_145_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12060_ _06047_ _06048_ _152_\[30\] VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__a21o_1
XFILLER_2_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11011_ net63 _04849_ _05147_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__a21o_1
XFILLER_2_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12962_ clknet_leaf_39_clk _00181_ VGND VGND VPWR VPWR _243_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11913_ _05906_ _05909_ _05904_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__o21ai_1
X_12893_ clknet_leaf_68_clk _00117_ VGND VGND VPWR VPWR _116_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11844_ _142_\[10\] _05853_ _05765_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__mux2_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11775_ _140_\[24\] _140_\[15\] VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__xnor2_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13514_ clknet_leaf_55_clk _00733_ VGND VGND VPWR VPWR _152_\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _170_\[15\] _04942_ _04922_ _04948_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__o211a_1
XFILLER_70_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10657_ _02476_ _04861_ _04900_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__a21boi_1
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13445_ clknet_leaf_127_clk _00664_ VGND VGND VPWR VPWR _164_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10588_ _173_\[4\] _176_\[4\] _01226_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__mux2_1
X_13376_ clknet_leaf_125_clk _00595_ VGND VGND VPWR VPWR _170_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12327_ _06195_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12258_ _06159_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__clkbuf_1
X_11209_ _05287_ _05288_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__nand2_1
XFILLER_122_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12189_ _01393_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__clkbuf_4
XFILLER_122_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06750_ _01321_ _01358_ _01403_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__or3_1
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06681_ _01372_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08420_ _02858_ _01801_ _02824_ _02859_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__o211a_1
XFILLER_91_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08351_ _228_\[11\] _02775_ _02753_ _02806_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__a211o_1
X_07302_ _182_\[5\] _01620_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__nor2_1
X_08282_ _228_\[26\] _02733_ _02723_ _02754_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__o211a_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07233_ _01790_ _01792_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__or2_1
XFILLER_118_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07164_ _01690_ _01726_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__xnor2_2
XFILLER_132_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07095_ _237_\[20\] VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__buf_6
XFILLER_133_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09805_ _04186_ _04190_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__and2_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07997_ _182_\[28\] _01698_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__nor2_1
X_09736_ _04124_ _04122_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__and2b_1
XFILLER_101_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06948_ _176_\[15\] _01531_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__or2_1
X_09667_ _03884_ _04058_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__or2_1
XFILLER_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06879_ _179_\[28\] _01302_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__or2_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _03045_ _03046_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__nor2_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09598_ _03989_ _03991_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__or2_1
XFILLER_91_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _02823_ _02787_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__xnor2_1
X_11560_ _05595_ _05597_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__xor2_1
XFILLER_11_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10511_ _179_\[13\] _04799_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__or2_1
XFILLER_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13230_ clknet_leaf_27_clk _00449_ VGND VGND VPWR VPWR _182_\[8\] sky130_fd_sc_hd__dfxtp_1
X_11491_ _05519_ _05530_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__or2_1
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10442_ _04685_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10373_ _179_\[5\] _04684_ _04686_ _04701_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__o211a_1
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13161_ clknet_leaf_109_clk _00380_ VGND VGND VPWR VPWR _225_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12112_ _140_\[17\] _142_\[17\] _06079_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__mux2_1
X_13092_ clknet_leaf_111_clk _00311_ VGND VGND VPWR VPWR _231_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12043_ _06030_ _06034_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__xor2_1
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12945_ clknet_leaf_21_clk _00164_ VGND VGND VPWR VPWR _246_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _118_\[29\] _120_\[29\] _06473_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__mux2_1
XFILLER_34_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _05835_ _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__nand2_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _142_\[3\] _05774_ _05765_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__mux2_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10709_ _01213_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__clkbuf_4
X_11689_ _116_\[28\] _05712_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__nand2_1
XFILLER_139_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13428_ clknet_leaf_123_clk _00647_ VGND VGND VPWR VPWR _164_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13359_ clknet_leaf_0_clk _00578_ VGND VGND VPWR VPWR _170_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07920_ _02424_ _02425_ _02456_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__a21oi_1
XFILLER_114_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07851_ _02364_ _02365_ _02388_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__and3_1
Xinput2 din[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
X_06802_ _246_\[7\] _01422_ _01425_ _01454_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__o211a_1
XFILLER_96_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07782_ _02303_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__inv_2
X_09521_ _185_\[0\] _03869_ _03379_ _03918_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__o211a_1
XFILLER_83_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06733_ _01400_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06664_ _01360_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__buf_4
XFILLER_101_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09452_ _03845_ _03855_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06595_ _099_ _01297_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__nand2_1
XFILLER_51_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08403_ net51 _02846_ _01353_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__mux2_1
X_09383_ _03746_ _03778_ _03787_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__nand3_1
XFILLER_52_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08334_ _228_\[7\] _02775_ _02753_ _02793_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__a211o_1
XFILLER_138_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08265_ _231_\[21\] _02730_ _02712_ _02742_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__a211o_1
X_07216_ _01774_ _01776_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__xnor2_1
X_08196_ _164_\[2\] _228_\[2\] _02687_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__mux2_1
XFILLER_118_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07147_ _182_\[0\] _237_\[0\] VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__nand2_2
XFILLER_145_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07078_ _173_\[16\] _01646_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__or2_1
XFILLER_114_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09719_ _03886_ _04103_ _04107_ _04108_ _04054_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__o2111a_1
XFILLER_90_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10991_ _164_\[29\] _05107_ _04865_ _05135_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__o211a_1
XFILLER_55_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12730_ _124_\[23\] _122_\[23\] _06401_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__mux2_1
XFILLER_15_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _126_\[22\] _124_\[22\] _06368_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__mux2_1
X_11612_ _118_\[23\] _118_\[27\] VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__xnor2_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12592_ _06334_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__clkbuf_1
X_11543_ _05582_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11474_ _05506_ _05511_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__or2_1
XFILLER_7_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13213_ clknet_leaf_41_clk _00432_ VGND VGND VPWR VPWR _185_\[23\] sky130_fd_sc_hd__dfxtp_4
X_10425_ _04712_ _04738_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__or2_1
XFILLER_109_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13144_ clknet_leaf_103_clk _00363_ VGND VGND VPWR VPWR _228_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10356_ _182_\[1\] _01217_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__or2_1
XFILLER_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _04637_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13075_ clknet_leaf_99_clk _00294_ VGND VGND VPWR VPWR _234_\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ _140_\[12\] _140_\[14\] VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__nand2_1
XFILLER_78_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13977_ clknet_leaf_91_clk _01196_ VGND VGND VPWR VPWR _118_\[25\] sky130_fd_sc_hd__dfxtp_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12928_ clknet_leaf_40_clk _00147_ VGND VGND VPWR VPWR _246_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _06474_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08050_ _02581_ _02582_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07001_ _01480_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__buf_2
XFILLER_115_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08952_ _170_\[16\] _02820_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__nand2_1
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07903_ _182_\[25\] _01687_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__nand2_1
X_08883_ _03244_ _03271_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__nand2_1
XFILLER_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07834_ _02334_ _02360_ _02372_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07765_ _02303_ _02306_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__xor2_1
X_09504_ _03874_ _01279_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__or2b_1
X_06716_ _01390_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__clkbuf_1
X_07696_ _01687_ _01642_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__xnor2_1
X_06647_ _01348_ VGND VGND VPWR VPWR _436_\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09435_ _03806_ _03809_ _03807_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__a21bo_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06578_ _01239_ _01286_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__nand2_1
X_09366_ _03771_ _03772_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__nand2_1
XANTENNA_40 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09297_ _01355_ _03696_ _03697_ _03705_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__a31o_1
X_08317_ _228_\[3\] _02771_ _02765_ _02780_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__o211a_1
XANTENNA_51 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _142_\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _01519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08248_ _01406_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__clkbuf_4
XFILLER_20_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10210_ _01233_ _04578_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__nand2_1
X_08179_ _231_\[29\] _02649_ _02679_ _02680_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__o211a_1
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11190_ _149_\[1\] _132_\[1\] VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__nand2_1
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10141_ _243_\[26\] _04409_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__or2_1
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10072_ _04411_ _04422_ _04446_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__or3_1
XFILLER_0_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13900_ clknet_leaf_97_clk _01119_ VGND VGND VPWR VPWR _122_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13831_ clknet_leaf_62_clk _01050_ VGND VGND VPWR VPWR _126_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13762_ clknet_leaf_63_clk _00981_ VGND VGND VPWR VPWR _130_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10974_ net51 _04853_ _05124_ _05117_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__o211a_1
XFILLER_46_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12713_ _124_\[15\] _122_\[15\] _06390_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__mux2_1
X_13693_ clknet_leaf_57_clk _00912_ VGND VGND VPWR VPWR _136_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12644_ _126_\[14\] _124_\[14\] _06357_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__mux2_1
XFILLER_31_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12575_ _128_\[13\] _126_\[13\] _06324_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__mux2_1
XFILLER_129_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11526_ _116_\[11\] _05566_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__nand2_1
XFILLER_144_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11457_ _116_\[4\] _05503_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__or2_1
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11388_ _05443_ _05444_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__nor2_1
X_10408_ _179_\[15\] _04721_ _04705_ _04726_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__o211a_1
XFILLER_140_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10339_ _179_\[29\] _04637_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__or2_1
XFILLER_3_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ clknet_leaf_106_clk _00346_ VGND VGND VPWR VPWR _228_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13058_ clknet_leaf_112_clk _00277_ VGND VGND VPWR VPWR _234_\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12009_ _01360_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__buf_6
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07550_ _02073_ _02074_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__and2b_1
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06501_ _01214_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__buf_6
X_07481_ _01924_ _01925_ _01964_ _02031_ _01943_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__o2111ai_4
XFILLER_62_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09220_ _03499_ _03534_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__nand2_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09151_ _03562_ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__and2_1
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09082_ _03479_ _03480_ _03496_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__o21ai_1
X_08102_ _01518_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__buf_4
XFILLER_135_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08033_ _182_\[30\] _01704_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__or2_1
XFILLER_116_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09984_ _04075_ _01284_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__nor2_1
XFILLER_115_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08935_ _03351_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__xnor2_1
X_08866_ _02074_ _03259_ _03286_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07817_ _182_\[23\] _01681_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__xor2_4
X_08797_ _02814_ _02776_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__xnor2_1
X_07748_ _02285_ _02287_ _02290_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__a21oi_1
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07679_ _02220_ _02223_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__xor2_2
XFILLER_53_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10690_ _173_\[5\] _04917_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__or2_1
X_09418_ _03821_ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__nor2_1
XFILLER_12_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09349_ _03718_ _03742_ _03755_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__a21oi_1
X_12360_ _06213_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11311_ _05368_ _05373_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__nand2_1
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12291_ _06176_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11242_ _01361_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__buf_4
XFILLER_134_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11173_ _05227_ _05257_ _05258_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__a21o_1
X_10124_ _04495_ _04496_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__or2_1
XFILLER_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10055_ _246_\[22\] _01315_ _04409_ _243_\[22\] _01497_ VGND VGND VPWR VPWR _04431_
+ sky130_fd_sc_hd__o221a_1
XFILLER_94_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13814_ clknet_leaf_94_clk _01033_ VGND VGND VPWR VPWR _128_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13745_ clknet_leaf_79_clk _00964_ VGND VGND VPWR VPWR _132_\[17\] sky130_fd_sc_hd__dfxtp_2
X_10957_ net45 _05110_ _05112_ _05086_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__a211o_1
X_13676_ clknet_leaf_77_clk _00895_ VGND VGND VPWR VPWR _136_\[12\] sky130_fd_sc_hd__dfxtp_1
X_12627_ _126_\[6\] _124_\[6\] _06346_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__mux2_1
X_10888_ _164_\[30\] _05048_ _05063_ _04998_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__o211a_1
XFILLER_145_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12558_ _128_\[5\] _126_\[5\] _06313_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__mux2_1
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12489_ _130_\[4\] _128_\[4\] _06280_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__mux2_1
X_11509_ _05549_ _05551_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__nand2_1
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06981_ _240_\[24\] _01565_ _01558_ _01584_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__o211a_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08720_ _01939_ _03108_ _03145_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__a21oi_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08651_ _03037_ _03039_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__and2b_1
XFILLER_39_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07602_ _01678_ _01632_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08582_ _01847_ _03011_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__xnor2_2
XFILLER_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07533_ _02081_ _02082_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__nand2_1
XFILLER_41_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07464_ _02014_ _02015_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__or2_1
X_09203_ _02383_ _03613_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__xor2_1
X_07395_ _01941_ _01944_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__nor2_1
XFILLER_50_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09134_ _02807_ _225_\[3\] VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09065_ _03453_ _03455_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__and2b_1
X_08016_ _02548_ _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09967_ _04345_ _04346_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__nand2_1
XFILLER_103_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08918_ _03336_ _03337_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__xnor2_2
X_09898_ _03905_ _04230_ _04280_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__a21o_1
XFILLER_94_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08849_ _170_\[13\] _02811_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__nand2_1
X_11860_ _152_\[12\] _05866_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__or2_1
XFILLER_45_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11791_ _152_\[6\] _05803_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__or2_1
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10811_ _04685_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__clkbuf_4
X_13530_ clknet_leaf_67_clk _00749_ VGND VGND VPWR VPWR _152_\[26\] sky130_fd_sc_hd__dfxtp_1
X_10742_ _167_\[19\] _04945_ _04960_ _04952_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__a211o_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13461_ clknet_leaf_123_clk _00680_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfxtp_4
X_10673_ _04888_ _04910_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__or2_1
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12412_ _06240_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__clkbuf_1
X_13392_ clknet_leaf_1_clk _00611_ VGND VGND VPWR VPWR _167_\[10\] sky130_fd_sc_hd__dfxtp_1
X_12343_ _06204_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12274_ _138_\[30\] _136_\[30\] _06167_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__mux2_1
X_11225_ _05289_ _05290_ _05295_ _05302_ _05294_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__o311a_1
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11156_ _158_\[16\] _01262_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10107_ _04161_ _04480_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__nor2_1
X_11087_ _05192_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10038_ _04078_ _04032_ _04383_ _04414_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__o31a_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13728_ clknet_leaf_66_clk _00947_ VGND VGND VPWR VPWR _132_\[0\] sky130_fd_sc_hd__dfxtp_1
X_11989_ _152_\[24\] _05983_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__or2_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13659_ clknet_leaf_56_clk _00878_ VGND VGND VPWR VPWR _138_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07180_ _01604_ _01742_ _01411_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__mux2_1
XFILLER_118_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09821_ _142_\[12\] _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__and2_1
XFILLER_113_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09752_ _04137_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__nor2_1
XFILLER_86_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06964_ _01568_ _01572_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__or2_1
XFILLER_55_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ _170_\[9\] _02797_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__nand2_1
X_09683_ _142_\[7\] _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06895_ _01353_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__clkbuf_8
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _02787_ _03032_ _02861_ _03062_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__a211o_1
XFILLER_82_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _02994_ _02995_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__and2_1
XFILLER_42_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07516_ _185_\[13\] _234_\[13\] VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__nand2_1
XFILLER_35_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08496_ _02904_ _02928_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__nand2_1
X_07447_ _01918_ _01921_ _01969_ _01999_ _01968_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__o311a_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07378_ _01931_ _01932_ _01930_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__a21o_1
XFILLER_6_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09117_ _03528_ _03530_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__xor2_1
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09048_ _03462_ _03463_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__xor2_2
XFILLER_123_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11010_ _164_\[5\] net68 _03030_ _04692_ _01417_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__a221o_1
XFILLER_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12961_ clknet_leaf_20_clk _00180_ VGND VGND VPWR VPWR _243_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12892_ clknet_leaf_68_clk _00116_ VGND VGND VPWR VPWR _116_\[1\] sky130_fd_sc_hd__dfxtp_1
X_11912_ _152_\[17\] _05914_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11843_ net2 _05851_ _05852_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__mux2_1
XFILLER_61_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11774_ _05789_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__clkbuf_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13513_ clknet_leaf_55_clk _00732_ VGND VGND VPWR VPWR _152_\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _173_\[15\] _04917_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__or2_1
XFILLER_14_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10656_ _176_\[26\] _04678_ _04627_ _173_\[26\] _02833_ VGND VGND VPWR VPWR _04900_
+ sky130_fd_sc_hd__o221a_1
X_13444_ clknet_leaf_128_clk _00663_ VGND VGND VPWR VPWR _164_\[30\] sky130_fd_sc_hd__dfxtp_1
X_10587_ _04686_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__buf_4
XFILLER_5_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13375_ clknet_leaf_127_clk _00594_ VGND VGND VPWR VPWR _170_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12326_ _136_\[23\] _134_\[23\] _06189_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__mux2_1
XFILLER_141_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12257_ _138_\[22\] _136_\[22\] _06156_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__mux2_1
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11208_ _149_\[4\] _132_\[4\] VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__nand2_1
X_12188_ _06122_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11139_ _158_\[12\] _01259_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__nand2_1
XFILLER_96_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06680_ _118_\[5\] _116_\[5\] _01370_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__mux2_1
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08350_ _02804_ _02791_ _02760_ _02805_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__o211a_1
XFILLER_24_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07301_ _01857_ _01858_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__nand2_1
X_08281_ _164_\[26\] _02736_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__or2_1
X_07232_ _01790_ _01792_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__nand2_1
XFILLER_20_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07163_ _01642_ _01626_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07094_ _01405_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__buf_2
XFILLER_132_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09804_ _04186_ _04190_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__nor2_1
XFILLER_101_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07996_ _02414_ _02528_ _02530_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__a21oi_2
X_09735_ _04122_ _04124_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__and2b_1
XFILLER_86_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06947_ _243_\[14\] _01536_ _01557_ _01560_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__a211o_1
XFILLER_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09666_ _03890_ _03896_ _03898_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__and3_1
XFILLER_39_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06878_ _01420_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__buf_2
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _228_\[6\] _231_\[6\] _02787_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__a21oi_2
X_09597_ _03989_ _03991_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__nand2_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _02960_ _02962_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__and2b_1
X_08479_ _02817_ _02781_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11490_ _05534_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__clkbuf_1
X_10510_ _01216_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__clkbuf_2
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10441_ _176_\[24\] _04725_ _04750_ _04728_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__a211o_1
XFILLER_109_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10372_ _182_\[5\] _04696_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__or2_1
X_13160_ clknet_leaf_109_clk _00379_ VGND VGND VPWR VPWR _225_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12111_ _06082_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__clkbuf_1
X_13091_ clknet_leaf_115_clk _00310_ VGND VGND VPWR VPWR _231_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12042_ _06032_ _06033_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__nor2_1
XFILLER_2_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12944_ clknet_leaf_39_clk _00163_ VGND VGND VPWR VPWR _246_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _06482_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _05836_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__inv_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11757_ net26 _05773_ _05742_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__mux2_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10708_ _167_\[10\] _04836_ _04935_ _04914_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__a211o_1
X_11688_ _118_\[3\] _05711_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10639_ _04681_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__clkbuf_2
X_13427_ clknet_leaf_123_clk _00646_ VGND VGND VPWR VPWR _164_\[13\] sky130_fd_sc_hd__dfxtp_1
X_13358_ clknet_leaf_11_clk _00577_ VGND VGND VPWR VPWR _170_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12309_ _136_\[15\] _134_\[15\] _06178_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__mux2_1
XFILLER_142_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13289_ clknet_leaf_24_clk _00508_ VGND VGND VPWR VPWR _176_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07850_ _02364_ _02365_ _02388_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06801_ _01444_ _01453_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__nand2_1
XFILLER_96_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07781_ _02310_ _02311_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__and2b_1
XFILLER_37_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09520_ _03870_ _03917_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__nand2_1
X_06732_ _118_\[29\] _116_\[29\] _01394_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__mux2_1
Xinput3 din[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
XFILLER_36_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06663_ _01321_ _01358_ _01359_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__or3b_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09451_ _03846_ _03854_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06594_ _158_\[21\] _01265_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__nor2_2
XFILLER_101_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08402_ _225_\[23\] VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__buf_6
X_09382_ _03746_ _03778_ _03787_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__a21o_1
XFILLER_24_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_125_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_125_clk sky130_fd_sc_hd__clkbuf_16
X_08333_ _02790_ _02791_ _02760_ _02792_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__o211a_1
X_08264_ _228_\[21\] _02733_ _02723_ _02741_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__o211a_1
X_07215_ _01749_ _01775_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__nor2_1
X_08195_ _231_\[1\] _02690_ _02664_ _02692_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__a211o_1
X_07146_ _01417_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__buf_4
XFILLER_133_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07077_ _237_\[16\] VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__buf_4
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09718_ _04002_ _01283_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__or2_1
XFILLER_75_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07979_ _243_\[28\] _240_\[28\] _01698_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__mux2_4
XFILLER_28_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10990_ _167_\[29\] _04867_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__or2_1
XFILLER_19_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09649_ _04038_ _04039_ _04041_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__and3_1
XFILLER_83_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12660_ _06370_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11611_ _05642_ _05643_ _149_\[19\] _05262_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12591_ _128_\[21\] _126_\[21\] _06324_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__mux2_1
XFILLER_11_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_116_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_116_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11542_ _149_\[12\] _05581_ _05533_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__mux2_1
XFILLER_137_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11473_ _05517_ _05518_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__nand2_1
XFILLER_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13212_ clknet_leaf_37_clk _00431_ VGND VGND VPWR VPWR _185_\[22\] sky130_fd_sc_hd__dfxtp_4
X_10424_ _179_\[20\] _182_\[20\] _04693_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__mux2_1
XFILLER_7_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13143_ clknet_leaf_119_clk _00362_ VGND VGND VPWR VPWR _228_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10355_ _176_\[0\] _04683_ _04688_ _01419_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__a211o_1
XFILLER_3_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _182_\[6\] _04634_ _04645_ _00105_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__o211a_1
XFILLER_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13074_ clknet_leaf_99_clk _00293_ VGND VGND VPWR VPWR _234_\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12025_ _140_\[12\] _140_\[14\] VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__or2_1
XFILLER_65_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13976_ clknet_leaf_91_clk _01195_ VGND VGND VPWR VPWR _118_\[24\] sky130_fd_sc_hd__dfxtp_2
X_12927_ clknet_leaf_30_clk _436_\[4\] _00104_ VGND VGND VPWR VPWR _392_\[4\] sky130_fd_sc_hd__dfstp_2
XFILLER_74_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12858_ _118_\[20\] _120_\[20\] _06473_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__mux2_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _140_\[25\] _140_\[27\] VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_107_clk sky130_fd_sc_hd__clkbuf_16
X_12789_ _122_\[19\] _120_\[19\] _06434_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__mux2_1
XFILLER_128_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07000_ _243_\[30\] _01548_ _01545_ _01597_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__o211a_1
XFILLER_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08951_ _170_\[16\] _02820_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__or2_1
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07902_ _02436_ _02438_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__or2_1
X_08882_ _03301_ _03302_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__and2b_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07833_ _02334_ _02360_ _02372_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__nor3_1
XFILLER_111_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07764_ _02304_ _02305_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__nand2_1
X_09503_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__clkbuf_4
X_06715_ _118_\[22\] _116_\[22\] _01381_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__mux2_1
X_07695_ _02215_ _02216_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__and2b_1
XFILLER_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06646_ _01338_ _01341_ _01343_ _01347_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__or4b_1
XFILLER_80_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09434_ _03837_ _03838_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__nand2_1
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06577_ _01244_ _01276_ _01285_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__and3_1
X_09365_ _170_\[28\] _02862_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__nand2_1
XFILLER_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_41 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09296_ _01427_ _03704_ _02002_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__a21o_1
X_08316_ _02749_ _02779_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__or2_1
XANTENNA_74 _142_\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _01635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08247_ _231_\[16\] _02706_ _02695_ _02729_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__o211a_1
XANTENNA_85 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08178_ _167_\[29\] _02652_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__or2_1
XFILLER_106_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07129_ _240_\[27\] _01649_ _01693_ _01697_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__a211o_1
X_10140_ _04497_ _04503_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10071_ _04411_ _04422_ _04446_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__o21ai_1
XFILLER_87_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13830_ clknet_leaf_61_clk _01049_ VGND VGND VPWR VPWR _126_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13761_ clknet_leaf_66_clk _00980_ VGND VGND VPWR VPWR _130_\[1\] sky130_fd_sc_hd__dfxtp_1
X_10973_ _05079_ _05123_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__or2_1
XFILLER_28_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12712_ _06397_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__clkbuf_1
X_13692_ clknet_leaf_57_clk _00911_ VGND VGND VPWR VPWR _136_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12643_ _06361_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12574_ _06325_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11525_ _118_\[18\] _05565_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11456_ _116_\[4\] _05503_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__nand2_1
XFILLER_124_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11387_ _149_\[27\] _132_\[27\] VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__and2_1
XFILLER_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10407_ _182_\[15\] _04696_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__or2_1
XFILLER_124_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10338_ _179_\[28\] _04658_ _04675_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__a21o_1
X_13126_ clknet_leaf_109_clk _00345_ VGND VGND VPWR VPWR _228_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13057_ clknet_leaf_15_clk _00276_ VGND VGND VPWR VPWR _234_\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12008_ net18 _05742_ _06001_ _06002_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__o22a_1
XFILLER_94_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10269_ _04633_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__clkbuf_4
XFILLER_93_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13959_ clknet_leaf_70_clk _01178_ VGND VGND VPWR VPWR _118_\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_81_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07480_ _01991_ _02021_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__nor2_1
X_06500_ _01213_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__buf_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09150_ _03545_ _03546_ _03561_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__or3_1
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09081_ _03493_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__xnor2_1
X_08101_ _01405_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__clkbuf_2
X_08032_ _182_\[30\] _01704_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__nand2_1
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09983_ _03901_ _04006_ _03873_ _03910_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__a31o_1
XFILLER_116_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08934_ _02127_ _03319_ _03352_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__a21oi_2
XFILLER_97_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08865_ _03256_ _03258_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__nor2_1
XFILLER_29_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08796_ _03197_ _02017_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__and2b_1
XFILLER_57_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07816_ _01678_ _01973_ _01886_ _02356_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__o211a_1
XFILLER_123_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07747_ _02288_ _02289_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__nand2_1
XFILLER_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07678_ _02166_ _02221_ _02222_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__o21ai_2
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06629_ _01323_ _01324_ _01325_ _01331_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__and4_1
XFILLER_52_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09417_ _03781_ _03785_ _03820_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__and3_1
XFILLER_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ _03753_ _03754_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__nand2_1
X_11310_ _05375_ _05376_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__or2b_1
X_09279_ _03685_ _03687_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12290_ _136_\[6\] _134_\[6\] _06167_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__mux2_1
XFILLER_113_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11241_ _05314_ _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__xor2_1
XFILLER_107_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11172_ net22 _05190_ _05192_ _158_\[20\] VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__a22o_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10123_ _142_\[25\] _04494_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__nor2_1
XFILLER_122_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10054_ _185_\[21\] _03870_ _03864_ _04430_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__o211a_1
XFILLER_102_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13813_ clknet_leaf_93_clk _01032_ VGND VGND VPWR VPWR _128_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13744_ clknet_leaf_79_clk _00963_ VGND VGND VPWR VPWR _132_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10956_ _164_\[18\] _05107_ _05094_ _05111_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__o211a_1
X_13675_ clknet_leaf_48_clk _00894_ VGND VGND VPWR VPWR _136_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10887_ _05028_ _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__or2_1
X_12626_ _06352_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12557_ _06316_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12488_ _06200_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__buf_6
X_11508_ _05550_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__inv_2
X_11439_ _116_\[1\] _05480_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__nand2_1
XFILLER_113_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ clknet_leaf_118_clk _00328_ VGND VGND VPWR VPWR _231_\[21\] sky130_fd_sc_hd__dfxtp_1
X_06980_ _176_\[24\] _01580_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__or2_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08650_ _01906_ _03077_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__xor2_2
XFILLER_39_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07601_ _02144_ _02147_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__nand2_1
XFILLER_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08581_ _03008_ _03010_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__xor2_4
XFILLER_47_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07532_ _182_\[13\] _01645_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__nand2_1
X_07463_ _01979_ _02007_ _02013_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__and3_1
XFILLER_62_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09202_ _185_\[24\] _03612_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__xnor2_1
X_07394_ _01407_ _01947_ _01948_ _00105_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__o211a_1
X_09133_ _03528_ _03530_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__and2_1
XFILLER_108_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09064_ _03450_ _03452_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__nor2_1
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08015_ _243_\[29\] _240_\[29\] _01701_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__mux2_4
XFILLER_118_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09966_ _04342_ _04344_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__or2_1
XFILLER_89_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09897_ _04078_ _04231_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__nand2_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08917_ _03301_ _03305_ _03302_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__o21ai_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08848_ _170_\[13\] _02811_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_96_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_73_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08779_ _228_\[11\] _231_\[11\] _03202_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__o21a_1
X_11790_ _152_\[6\] _05803_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__nand2_1
X_10810_ _164_\[7\] _04983_ _05008_ _04998_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__o211a_1
XFILLER_53_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10741_ _170_\[19\] _04942_ _04958_ _04959_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__o211a_1
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13460_ clknet_leaf_114_clk _00679_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_2
XFILLER_139_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12411_ _132_\[31\] _134_\[31\] _06230_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__mux2_1
X_10672_ _170_\[0\] _173_\[0\] _04830_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_20_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
X_13391_ clknet_leaf_2_clk _00610_ VGND VGND VPWR VPWR _167_\[9\] sky130_fd_sc_hd__dfxtp_2
X_12342_ _136_\[30\] _134_\[30\] _06201_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__mux2_1
XFILLER_5_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12273_ _01393_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__clkbuf_4
XFILLER_5_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11224_ _149_\[4\] _132_\[4\] _05293_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__nand3_1
XFILLER_5_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11155_ _05245_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10106_ _04436_ _04479_ _03906_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__a21oi_1
X_11086_ _05190_ _05191_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__nor2_4
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10037_ _01244_ _03878_ _03976_ _03897_ _01237_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__a2111o_1
XFILLER_76_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_87_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_91_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11988_ _152_\[24\] _05983_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__nand2_1
XFILLER_63_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13727_ clknet_leaf_58_clk _00946_ VGND VGND VPWR VPWR _134_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10939_ _164_\[13\] _05059_ _05094_ _05099_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__o211a_1
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13658_ clknet_leaf_56_clk _00877_ VGND VGND VPWR VPWR _138_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13589_ clknet_leaf_50_clk _00808_ VGND VGND VPWR VPWR _142_\[21\] sky130_fd_sc_hd__dfxtp_1
X_12609_ _06343_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_31_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09820_ _246_\[12\] _01314_ _03914_ _243_\[12\] _01466_ VGND VGND VPWR VPWR _04206_
+ sky130_fd_sc_hd__o221a_1
XFILLER_140_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09751_ _04103_ _04010_ _04138_ _04139_ _04078_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__o221a_1
XFILLER_101_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06963_ _176_\[19\] _240_\[19\] _01569_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__mux2_1
XFILLER_140_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_78_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_16
X_08702_ _170_\[9\] _02797_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__or2_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09682_ _246_\[7\] _01314_ _03914_ _243_\[7\] _01452_ VGND VGND VPWR VPWR _04073_
+ sky130_fd_sc_hd__o221a_1
X_06894_ _246_\[31\] _01485_ _01481_ _01522_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__o211a_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08633_ _02380_ _03053_ _03061_ _02202_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__o211a_1
XFILLER_27_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _02978_ _02979_ _02993_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__or3_1
XFILLER_23_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07515_ _185_\[13\] _234_\[13\] VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__or2_1
X_08495_ _02925_ _02927_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__xor2_2
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07446_ _182_\[8\] _01629_ _01967_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__nand3_1
XFILLER_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07377_ _01930_ _01931_ _01932_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__nand3_1
XFILLER_10_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09116_ _228_\[21\] _231_\[21\] _03529_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__o21a_1
X_09047_ _03436_ _03437_ _03435_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09949_ _04329_ _04311_ _04308_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__and3b_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_69_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12960_ clknet_leaf_43_clk _00179_ VGND VGND VPWR VPWR _243_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11911_ _140_\[27\] _05913_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__xnor2_2
X_12891_ clknet_leaf_68_clk _00115_ VGND VGND VPWR VPWR _116_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11842_ _01358_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__buf_4
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11773_ _142_\[4\] _05788_ _05765_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__mux2_1
X_13512_ clknet_leaf_55_clk _00731_ VGND VGND VPWR VPWR _152_\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10724_ _167_\[14\] _04945_ _04947_ _04914_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__a211o_1
X_10655_ _04861_ _04898_ _04899_ _04891_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__o211a_1
XFILLER_9_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13443_ clknet_leaf_122_clk _00662_ VGND VGND VPWR VPWR _164_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13374_ clknet_leaf_126_clk _00593_ VGND VGND VPWR VPWR _170_\[24\] sky130_fd_sc_hd__dfxtp_1
X_12325_ _06194_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__clkbuf_1
X_10586_ _173_\[3\] _04849_ _04852_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__a21o_1
XFILLER_142_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12256_ _06158_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__clkbuf_1
X_11207_ _149_\[4\] _132_\[4\] VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__or2_1
X_12187_ _140_\[21\] _138_\[21\] _06112_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__mux2_1
XFILLER_79_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11138_ _05227_ _05231_ _05232_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__a21o_1
XFILLER_95_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11069_ _164_\[28\] _03774_ _04636_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_0_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_91_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07300_ _182_\[6\] _01623_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__nand2_1
XFILLER_44_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08280_ _02711_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07231_ _01759_ _01760_ _01791_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__o21bai_1
X_07162_ _01725_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07093_ _240_\[19\] _01660_ _01653_ _01669_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__o211a_1
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09803_ _04188_ _04189_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__or2_1
XFILLER_115_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07995_ _02472_ _02479_ _02480_ _02529_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__o211ai_1
X_09734_ _04067_ _04066_ _04068_ _04095_ _04123_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__o41ai_2
XFILLER_101_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06946_ _240_\[14\] _01526_ _01558_ _01559_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__o211a_1
X_09665_ _03884_ _03901_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__nand2_1
XFILLER_95_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06877_ _01435_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__clkbuf_4
XFILLER_55_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08616_ _228_\[6\] _231_\[6\] VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__nor2_1
X_09596_ _03920_ _03942_ _03990_ _03968_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__a31o_1
XFILLER_131_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08547_ _02957_ _02959_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__nor2_1
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08478_ _01755_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__inv_2
X_07429_ _01954_ _01975_ _01981_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__a21o_1
XFILLER_7_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10440_ _179_\[24\] _04721_ _04705_ _04749_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__o211a_1
XFILLER_7_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10371_ _176_\[4\] _04691_ _04700_ _04677_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__o211a_1
XFILLER_40_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12110_ _140_\[16\] _142_\[16\] _06079_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__mux2_1
XFILLER_2_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13090_ clknet_leaf_115_clk _00309_ VGND VGND VPWR VPWR _231_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12041_ _152_\[28\] _06031_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__nor2_1
XFILLER_105_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12943_ clknet_leaf_21_clk _00162_ VGND VGND VPWR VPWR _246_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _118_\[28\] _120_\[28\] _06473_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__mux2_1
XFILLER_61_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _152_\[9\] _05834_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__nor2_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _05771_ _05772_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__xnor2_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10707_ _170_\[10\] _04833_ _04922_ _04934_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__o211a_1
X_11687_ _118_\[14\] _118_\[31\] VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__xnor2_1
X_13426_ clknet_leaf_113_clk _00645_ VGND VGND VPWR VPWR _164_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10638_ _04861_ _04886_ _04887_ _04823_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__o211a_1
XFILLER_142_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10569_ _173_\[29\] _04818_ _04841_ _04823_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__o211a_1
X_13357_ clknet_leaf_0_clk _00576_ VGND VGND VPWR VPWR _170_\[7\] sky130_fd_sc_hd__dfxtp_1
X_12308_ _06185_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__clkbuf_1
X_13288_ clknet_leaf_24_clk _00507_ VGND VGND VPWR VPWR _176_\[2\] sky130_fd_sc_hd__dfxtp_2
X_12239_ _06149_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06800_ _243_\[7\] _01428_ _01452_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__o21ai_1
X_07780_ _01675_ _01973_ _01886_ _02321_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__o211a_1
XFILLER_37_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 din[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
X_06731_ _01399_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09450_ _03851_ _03853_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__xnor2_1
X_06662_ _01302_ _01253_ _01309_ _01324_ net35 VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__a41o_1
XFILLER_64_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08401_ _01799_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__buf_4
XFILLER_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06593_ _01284_ _01296_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09381_ _03785_ _03786_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__nand2_1
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08332_ net65 _02736_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__or2_1
XFILLER_138_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08263_ _164_\[21\] _02736_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__or2_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07214_ _01711_ _01739_ _01747_ _01745_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__o211a_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08194_ _228_\[1\] _02649_ _02679_ _02691_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__o211a_1
XFILLER_20_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07145_ _240_\[31\] _01649_ _01693_ _01709_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__a211o_1
XFILLER_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07076_ _240_\[15\] _01601_ _01653_ _01656_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__o211a_1
XFILLER_133_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07978_ _02511_ _02512_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__or2_1
X_09717_ _01242_ _03890_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__nand2_2
X_06929_ _243_\[9\] _01485_ _01545_ _01547_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__o211a_1
XFILLER_87_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09648_ _03996_ _04018_ _04040_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__o21ai_1
XFILLER_55_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09579_ _246_\[3\] _01313_ _03914_ _243_\[3\] _01440_ VGND VGND VPWR VPWR _03974_
+ sky130_fd_sc_hd__o221a_2
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11610_ _05629_ _05634_ _05641_ _05352_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__a31o_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12590_ _06333_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11541_ _05578_ _05580_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__xor2_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11472_ _116_\[6\] _05516_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__or2_1
XFILLER_7_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13211_ clknet_leaf_41_clk _00430_ VGND VGND VPWR VPWR _185_\[21\] sky130_fd_sc_hd__dfxtp_2
X_10423_ _176_\[19\] _04735_ _04737_ _04677_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__o211a_1
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10354_ _179_\[0\] _04684_ _04686_ _04687_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__o211a_1
X_13142_ clknet_leaf_120_clk _00361_ VGND VGND VPWR VPWR _228_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10285_ _179_\[6\] _04638_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__or2_1
XFILLER_3_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13073_ clknet_leaf_99_clk _00292_ VGND VGND VPWR VPWR _234_\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12024_ _06017_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13975_ clknet_leaf_92_clk _01194_ VGND VGND VPWR VPWR _118_\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_19_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12926_ clknet_leaf_31_clk _436_\[3\] _00103_ VGND VGND VPWR VPWR _392_\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12857_ _06004_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__clkbuf_4
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11808_ _142_\[7\] _05279_ _05820_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__o21a_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12788_ _06437_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__clkbuf_1
X_11739_ _140_\[19\] _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13409_ clknet_leaf_126_clk _00628_ VGND VGND VPWR VPWR _167_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08950_ _03359_ _03368_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07901_ _02436_ _02438_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__nand2_1
X_08881_ _170_\[14\] _02814_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__nand2_1
XFILLER_111_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07832_ _02370_ _02371_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09502_ _01279_ _03874_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__or2b_1
XFILLER_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07763_ _185_\[21\] _234_\[21\] VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__nand2_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06714_ _01389_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__clkbuf_1
X_07694_ _02220_ _02223_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__nand2_1
XFILLER_37_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06645_ _190_\[3\] _01222_ _01345_ _01207_ _01346_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__o221a_1
XFILLER_64_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09433_ _170_\[30\] _02868_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__or2_1
XFILLER_24_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09364_ _170_\[28\] _02862_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__or2_1
XFILLER_13_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06576_ _01278_ _01281_ _01284_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__and3_1
XFILLER_12_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08315_ net61 _225_\[3\] _02750_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__mux2_1
XFILLER_138_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_31 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 _173_\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09295_ _03700_ _03703_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_64 _02001_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 _170_\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08246_ _02686_ _02728_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__or2_1
XFILLER_20_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_86 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08177_ _01420_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__clkbuf_4
XFILLER_119_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07128_ _01694_ _01639_ _01695_ _01696_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__o211a_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07059_ _173_\[12\] _01642_ _01617_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10070_ _04444_ _04445_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__and2b_1
XFILLER_88_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13760_ clknet_leaf_65_clk _00979_ VGND VGND VPWR VPWR _130_\[0\] sky130_fd_sc_hd__dfxtp_1
X_10972_ _164_\[23\] _167_\[23\] _01214_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__mux2_1
X_13691_ clknet_leaf_57_clk _00910_ VGND VGND VPWR VPWR _136_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12711_ _124_\[14\] _122_\[14\] _06390_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__mux2_1
XFILLER_102_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12642_ _126_\[13\] _124_\[13\] _06357_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__mux2_1
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12573_ _128_\[12\] _126_\[12\] _06324_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__mux2_1
XFILLER_23_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11524_ _118_\[14\] _118_\[29\] VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11455_ _118_\[7\] _05502_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10406_ _04724_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__buf_2
XFILLER_124_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11386_ _149_\[27\] _132_\[27\] VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__nor2_1
X_10337_ _182_\[28\] _04654_ _04671_ _01710_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__a31o_1
X_13125_ clknet_leaf_111_clk _00344_ VGND VGND VPWR VPWR _228_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10268_ _04626_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__buf_4
X_13056_ clknet_leaf_13_clk _00275_ VGND VGND VPWR VPWR _234_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12007_ _05999_ _06000_ _05785_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__o21ai_1
XFILLER_78_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10199_ _04554_ _04555_ _04556_ _04531_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__a22o_1
XFILLER_93_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13958_ clknet_leaf_72_clk _01177_ VGND VGND VPWR VPWR _118_\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_81_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12909_ clknet_leaf_86_clk _00133_ VGND VGND VPWR VPWR _116_\[18\] sky130_fd_sc_hd__dfxtp_1
X_13889_ clknet_leaf_69_clk _01108_ VGND VGND VPWR VPWR _122_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08100_ _234_\[6\] _02448_ _02419_ _02624_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__o211a_1
X_09080_ _228_\[20\] _231_\[20\] _03494_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__o21a_1
X_08031_ _01406_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__clkbuf_4
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09982_ _04075_ _03928_ _04078_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__o21ai_1
XFILLER_115_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08933_ _03316_ _03318_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__nor2_1
XFILLER_123_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08864_ _02097_ _03284_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08795_ _03194_ _03196_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__nor2_1
X_07815_ _02346_ _02347_ _02354_ _02355_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__a211o_1
XFILLER_29_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07746_ _182_\[20\] _01671_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__nand2_1
XFILLER_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07677_ _02198_ _02194_ _02196_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__a21o_1
XFILLER_53_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09416_ _03781_ _03785_ _03820_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__a21oi_1
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06628_ _01326_ _01330_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__nor2_1
XFILLER_52_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06559_ _01267_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__buf_4
X_09347_ _02514_ _03752_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__or2_1
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09278_ _228_\[26\] _231_\[26\] _03686_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__o21a_1
XFILLER_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08229_ _164_\[11\] _228_\[11\] _02687_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__mux2_1
XFILLER_119_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11240_ _05301_ _05303_ _05308_ _05315_ _05307_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__o311a_1
XFILLER_134_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11171_ _01265_ _05256_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__nand2_1
XFILLER_134_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10122_ _142_\[25\] _04494_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__and2_1
X_10053_ _04427_ _04428_ _04429_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__a21o_1
XFILLER_94_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13812_ clknet_leaf_94_clk _01031_ VGND VGND VPWR VPWR _128_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13743_ clknet_leaf_79_clk _00962_ VGND VGND VPWR VPWR _132_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10955_ _167_\[18\] _05089_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__or2_1
X_13674_ clknet_leaf_48_clk _00893_ VGND VGND VPWR VPWR _136_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10886_ _167_\[30\] _170_\[30\] _04995_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__mux2_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12625_ _126_\[5\] _124_\[5\] _06346_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__mux2_1
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12556_ _128_\[4\] _126_\[4\] _06313_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__mux2_1
XFILLER_12_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11507_ _116_\[9\] _05548_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__nor2_1
X_12487_ _06279_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__clkbuf_1
X_11438_ _05486_ _05487_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__or2b_1
XFILLER_140_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11369_ _05426_ _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__nand2_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13108_ clknet_leaf_104_clk _00327_ VGND VGND VPWR VPWR _231_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13039_ clknet_4_9_0_clk _00258_ VGND VGND VPWR VPWR _237_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07600_ _02032_ _02034_ _02145_ _02146_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__a211o_1
X_08580_ _01835_ _02982_ _03009_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__o21a_1
XFILLER_82_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07531_ _182_\[13\] _01645_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__or2_1
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07462_ _01979_ _02007_ _02013_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07393_ _01480_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__buf_4
XFILLER_22_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09201_ _02855_ _03611_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__xnor2_1
X_09132_ _03514_ _03515_ _03527_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__a21oi_1
XFILLER_118_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09063_ _03476_ _03477_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__nor2_1
X_08014_ _02546_ _02547_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__or2_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09965_ _04342_ _04344_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__nand2_1
X_09896_ _04011_ _04278_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__or2b_1
XFILLER_57_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08916_ _03334_ _03335_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__nor2_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08847_ _03251_ _03241_ _03267_ _01408_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__a31o_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08778_ _228_\[11\] _231_\[11\] _02804_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__a21o_1
X_07729_ _02270_ _02271_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10740_ _173_\[19\] _04953_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__or2_1
X_10671_ _04907_ _04909_ _03866_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__a21oi_1
X_12410_ _06239_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13390_ clknet_leaf_12_clk _00609_ VGND VGND VPWR VPWR _167_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12341_ _06203_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__clkbuf_1
X_12272_ _06166_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11223_ _05299_ _05300_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__nand2_1
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11154_ _05243_ _05244_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__or2_1
XFILLER_1_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10105_ _04320_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__inv_2
X_11085_ net35 _01248_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__nor2_4
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10036_ _04411_ _04412_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__or2_1
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11987_ _140_\[11\] _140_\[9\] VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__xor2_1
XFILLER_63_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13726_ clknet_leaf_57_clk _00945_ VGND VGND VPWR VPWR _134_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10938_ _167_\[13\] _05089_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__or2_1
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13657_ clknet_leaf_56_clk _00876_ VGND VGND VPWR VPWR _138_\[25\] sky130_fd_sc_hd__dfxtp_1
X_10869_ _164_\[24\] _05048_ _05050_ _04998_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__o211a_1
XFILLER_31_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13588_ clknet_leaf_46_clk _00807_ VGND VGND VPWR VPWR _142_\[20\] sky130_fd_sc_hd__dfxtp_1
X_12608_ _128_\[29\] _126_\[29\] _06335_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__mux2_1
XFILLER_8_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12539_ _130_\[28\] _128_\[28\] _06302_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__mux2_1
XFILLER_144_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09750_ _01242_ _03873_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__nand2_1
XFILLER_100_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06962_ _243_\[18\] _01548_ _01545_ _01571_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__o211a_1
X_09681_ _04049_ _04062_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__and2b_1
X_08701_ _02794_ _02845_ _02834_ _03127_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__o211a_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06893_ _243_\[31\] _01520_ _01495_ _01521_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__a211o_1
XFILLER_66_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08632_ _02404_ _03060_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__nand2_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08563_ _02978_ _02979_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__o21ai_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07514_ _02063_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__inv_2
X_08494_ _02900_ _02902_ _02926_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__a21o_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07445_ _01996_ _01997_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__nand2_1
XFILLER_50_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07376_ _185_\[8\] _234_\[8\] VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__nand2_1
XFILLER_10_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09115_ _228_\[21\] _231_\[21\] _02839_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__a21o_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09046_ _170_\[19\] _02830_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__xor2_2
XFILLER_145_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09948_ _04327_ _04328_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__xnor2_1
X_09879_ _04252_ _04261_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__nor2_1
XFILLER_58_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11910_ _140_\[2\] _140_\[4\] VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__xnor2_2
X_12890_ _06491_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11841_ _05847_ _05850_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__xor2_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11772_ net27 _05776_ _05784_ _05787_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__a22o_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13511_ clknet_leaf_60_clk _00730_ VGND VGND VPWR VPWR _152_\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10723_ _170_\[14\] _04942_ _04922_ _04946_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__o211a_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10654_ _02445_ _04724_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__nand2_1
XFILLER_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13442_ clknet_leaf_126_clk _00661_ VGND VGND VPWR VPWR _164_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10585_ _176_\[3\] net68 _01777_ _04692_ _02711_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__a221o_1
X_13373_ clknet_leaf_129_clk _00592_ VGND VGND VPWR VPWR _170_\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_126_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12324_ _136_\[22\] _134_\[22\] _06189_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__mux2_1
XFILLER_5_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12255_ _138_\[21\] _136_\[21\] _06156_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__mux2_1
X_11206_ _05279_ _05284_ _05285_ _05286_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__a31o_1
XFILLER_123_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12186_ _06121_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11137_ net13 _05202_ _05193_ _158_\[11\] VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__a22o_1
XFILLER_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11068_ net55 _04848_ _05182_ _01436_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__a211o_1
XFILLER_37_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10019_ _04310_ _04329_ _04396_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__or3b_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13709_ clknet_leaf_78_clk _00928_ VGND VGND VPWR VPWR _134_\[13\] sky130_fd_sc_hd__dfxtp_1
X_07230_ _01761_ _01762_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__and2b_1
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07161_ _01710_ _01724_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__or2_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07092_ _01615_ _01668_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__or2_1
XFILLER_133_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09802_ _142_\[11\] _04187_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__nor2_1
XFILLER_115_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07994_ _02406_ _02441_ _02527_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__a21o_1
X_09733_ _04096_ _04093_ _04094_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__a21bo_1
XFILLER_86_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06945_ _176_\[14\] _01531_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__or2_1
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09664_ _01284_ _04055_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__nand2_1
XFILLER_131_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06876_ _246_\[27\] _01496_ _01460_ _01508_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__a211o_1
XFILLER_67_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09595_ _03948_ _03949_ _03967_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__or3_1
X_08615_ _03041_ _03043_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__xnor2_2
XFILLER_55_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08546_ _02974_ _02976_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__xnor2_2
X_08477_ _02910_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__clkbuf_1
X_07428_ _01977_ _01980_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__xor2_1
XFILLER_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07359_ _01626_ _01660_ _01886_ _01915_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__o211a_1
XFILLER_7_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10370_ _04692_ _04699_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__or2_1
X_09029_ _185_\[19\] _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__xnor2_1
X_12040_ _152_\[28\] _06031_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__and2_1
XFILLER_120_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12942_ clknet_leaf_39_clk _00161_ VGND VGND VPWR VPWR _246_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12873_ _06481_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _152_\[9\] _05834_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__nand2_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _05759_ _05762_ _05758_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__a21bo_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _173_\[10\] _04917_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__or2_1
XFILLER_41_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11686_ _05710_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__clkbuf_1
X_13425_ clknet_leaf_1_clk _00644_ VGND VGND VPWR VPWR _164_\[11\] sky130_fd_sc_hd__dfxtp_2
X_10637_ _02293_ _04724_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__nand2_1
XFILLER_10_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10568_ _04809_ _04840_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__or2_1
X_13356_ clknet_leaf_3_clk _00575_ VGND VGND VPWR VPWR _170_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12307_ _136_\[14\] _134_\[14\] _06178_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__mux2_1
X_10499_ _04766_ _04791_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__or2_1
X_13287_ clknet_leaf_24_clk _00506_ VGND VGND VPWR VPWR _176_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12238_ _138_\[13\] _136_\[13\] _06145_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__mux2_1
XFILLER_111_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12169_ _140_\[12\] _138_\[12\] _06112_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__mux2_1
XFILLER_68_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput5 din[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
X_06730_ _118_\[28\] _116_\[28\] _01394_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__mux2_1
XFILLER_77_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06661_ _01273_ _01247_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__nor2_4
XFILLER_37_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08400_ _228_\[22\] _02838_ _02810_ _02844_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__a211o_1
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06592_ _01295_ _01253_ _01275_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__o21a_1
XFILLER_91_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09380_ _02540_ _03784_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__or2_1
XFILLER_36_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08331_ _01437_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__buf_2
X_08262_ _231_\[20\] _02706_ _02695_ _02740_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__o211a_1
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07213_ _01772_ _01773_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__or2b_1
XFILLER_20_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08193_ _164_\[1\] _02652_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__or2_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07144_ _01707_ _01639_ _01695_ _01708_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__o211a_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07075_ _01615_ _01655_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__or2_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07977_ _02488_ _02489_ _02510_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__and3_1
X_09716_ _01236_ _04102_ _04104_ _04105_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__a31o_1
X_06928_ _01448_ _01546_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__or2_1
XFILLER_74_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09647_ _04015_ _04017_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__or2b_1
X_06859_ _179_\[22\] _01301_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__or2_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09578_ _142_\[2\] _03965_ _03966_ _03964_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08529_ _228_\[3\] _231_\[3\] _225_\[3\] VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__a21o_1
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11540_ _05560_ _05562_ _05570_ _05579_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__o31a_1
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11471_ _116_\[6\] _05516_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__nand2_1
XFILLER_51_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13210_ clknet_leaf_41_clk _00429_ VGND VGND VPWR VPWR _185_\[20\] sky130_fd_sc_hd__dfxtp_4
X_10422_ _04712_ _04736_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__or2_1
XFILLER_137_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10353_ _182_\[0\] _01217_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__or2_1
X_13141_ clknet_leaf_118_clk _00360_ VGND VGND VPWR VPWR _228_\[21\] sky130_fd_sc_hd__dfxtp_1
X_13072_ clknet_leaf_99_clk _00291_ VGND VGND VPWR VPWR _234_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12023_ _142_\[26\] _06016_ _06005_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__mux2_1
X_10284_ _182_\[5\] _04634_ _04644_ _00105_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__o211a_1
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13974_ clknet_leaf_91_clk _01193_ VGND VGND VPWR VPWR _118_\[22\] sky130_fd_sc_hd__dfxtp_2
X_12925_ clknet_leaf_32_clk _436_\[2\] _00102_ VGND VGND VPWR VPWR _392_\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12856_ _06472_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__clkbuf_1
X_11807_ net30 _05776_ _05818_ _05819_ _01368_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__a221o_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _122_\[18\] _120_\[18\] _06434_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__mux2_1
X_11738_ _140_\[21\] _140_\[12\] VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11669_ _116_\[26\] _05693_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__or2_1
X_13408_ clknet_leaf_126_clk _00627_ VGND VGND VPWR VPWR _167_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13339_ clknet_leaf_0_clk _00558_ VGND VGND VPWR VPWR _173_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07900_ _02437_ _02402_ _02394_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__o21ai_1
X_08880_ _170_\[14\] _02814_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__nor2_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07831_ _243_\[23\] _240_\[23\] _01681_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__mux2_4
XFILLER_96_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09501_ _01241_ _03896_ _03898_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__and3_1
XFILLER_65_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07762_ _185_\[21\] _234_\[21\] VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__or2_1
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07693_ _02235_ _02236_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__xnor2_4
X_06713_ _118_\[21\] _116_\[21\] _01381_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__mux2_1
X_06644_ _01310_ _01324_ _01295_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__mux2_1
X_09432_ _170_\[30\] _02868_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__nand2_1
X_06575_ _01283_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__clkbuf_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09363_ _03701_ _03665_ _03767_ _03769_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__a31o_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08314_ _228_\[2\] _02775_ _02753_ _02778_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__a211o_1
XFILLER_33_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_32 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _179_\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 _05079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09294_ _03701_ _03664_ _03702_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__a21o_1
XANTENNA_65 _02001_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08245_ _164_\[16\] _228_\[16\] _02687_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__mux2_1
XANTENNA_43 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_76 _173_\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08176_ _234_\[28\] _02659_ _02636_ _02678_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__o211a_1
XFILLER_20_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_87 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07127_ _173_\[27\] _01646_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__or2_1
XFILLER_137_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07058_ _237_\[12\] VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__buf_4
XFILLER_133_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10971_ net50 _05110_ _05121_ _05122_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__a211o_1
X_13690_ clknet_leaf_56_clk _00909_ VGND VGND VPWR VPWR _136_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12710_ _06396_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12641_ _06360_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__clkbuf_1
X_12572_ _06200_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__clkbuf_4
XFILLER_11_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11523_ _05564_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11454_ _118_\[22\] _118_\[11\] VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10405_ _04681_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__buf_4
XFILLER_137_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11385_ _05441_ _05437_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__and2_1
X_10336_ _179_\[27\] _04658_ _04674_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__a21o_1
X_13124_ clknet_leaf_112_clk _00343_ VGND VGND VPWR VPWR _228_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10267_ _179_\[0\] _04629_ _04632_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__a21o_1
Xclkbuf_4_9_0_clk clknet_3_4_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_13055_ clknet_leaf_85_clk _00274_ VGND VGND VPWR VPWR _237_\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12006_ _05999_ _06000_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__and2_1
XFILLER_39_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10198_ _04554_ _04555_ _04556_ _04531_ _04567_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__a221oi_4
XFILLER_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13957_ clknet_leaf_71_clk _01176_ VGND VGND VPWR VPWR _118_\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12908_ clknet_leaf_86_clk _00132_ VGND VGND VPWR VPWR _116_\[17\] sky130_fd_sc_hd__dfxtp_1
X_13888_ clknet_leaf_69_clk _01107_ VGND VGND VPWR VPWR _122_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12839_ _118_\[11\] _120_\[11\] _06462_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__mux2_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08030_ _01701_ _02448_ _02419_ _02563_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__o211a_1
Xinput30 din[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
XFILLER_128_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09981_ _03878_ _04132_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__and2_1
XFILLER_115_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08932_ _03349_ _03350_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__or2_1
XFILLER_85_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08863_ _03281_ _03283_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__xor2_1
XFILLER_123_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08794_ _02804_ _02845_ _02834_ _03217_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__o211a_1
X_07814_ _01405_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__buf_4
XFILLER_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07745_ _182_\[20\] _01671_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__or2_1
XFILLER_53_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07676_ _02197_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__inv_2
XFILLER_53_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09415_ _03814_ _03819_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06627_ net35 _01327_ _01328_ _01329_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__or4_1
X_06558_ _392_\[0\] _392_\[4\] _392_\[1\] VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__or3b_1
X_09346_ _02514_ _03752_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__nand2_1
X_09277_ _228_\[26\] _231_\[26\] _02855_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__a21o_1
XFILLER_21_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08228_ _231_\[10\] _02706_ _02695_ _02716_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__o211a_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08159_ _167_\[23\] _231_\[23\] _02626_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__mux2_1
X_11170_ _158_\[19\] _01264_ _158_\[20\] VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__o21ai_1
XFILLER_134_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10121_ _246_\[25\] _01316_ _04409_ _243_\[25\] _01503_ VGND VGND VPWR VPWR _04494_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10052_ _04427_ _04428_ _03867_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13811_ clknet_leaf_95_clk _01030_ VGND VGND VPWR VPWR _128_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13742_ clknet_leaf_78_clk _00961_ VGND VGND VPWR VPWR _132_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10954_ _04682_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13673_ clknet_leaf_54_clk _00892_ VGND VGND VPWR VPWR _136_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10885_ _164_\[29\] _05025_ _05061_ _05035_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__a211o_1
X_12624_ _06351_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__clkbuf_1
X_12555_ _06315_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11506_ _116_\[9\] _05548_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__nand2_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12486_ _130_\[3\] _128_\[3\] _06269_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__mux2_1
XFILLER_8_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11437_ _116_\[2\] _05485_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__or2_1
XFILLER_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11368_ _149_\[25\] _132_\[25\] VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__or2_1
XFILLER_113_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10319_ _182_\[19\] _04663_ _04665_ _04649_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__o211a_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ clknet_leaf_118_clk _00326_ VGND VGND VPWR VPWR _231_\[19\] sky130_fd_sc_hd__dfxtp_1
X_11299_ _05367_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13038_ clknet_4_9_0_clk _00257_ VGND VGND VPWR VPWR _237_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07530_ _02078_ _02079_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07461_ _02009_ _02012_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__xor2_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07392_ _01629_ _01412_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__or2_1
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09200_ _02814_ _02784_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__xnor2_1
X_09131_ _03541_ _03543_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__xnor2_2
X_09062_ _03475_ _03469_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__and2b_1
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08013_ _02544_ _02545_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__and2_1
XFILLER_116_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09964_ _142_\[17\] _04325_ _04343_ _04324_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__a22o_1
X_09895_ _01242_ _04082_ _03936_ _01236_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__o31a_1
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08915_ _170_\[15\] _02817_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__and2_1
XFILLER_85_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _03251_ _03241_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__a21oi_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08777_ _03198_ _03200_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07728_ _243_\[20\] _240_\[20\] _01671_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__mux2_4
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07659_ _02191_ _02192_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__and2b_1
XFILLER_13_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10670_ _02606_ _04872_ _04637_ _04908_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__a211o_1
XFILLER_41_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09329_ _03731_ _03732_ _03736_ _01439_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__o211a_1
XFILLER_138_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12340_ _136_\[29\] _134_\[29\] _06201_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__mux2_1
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12271_ _138_\[29\] _136_\[29\] _06156_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__mux2_1
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11222_ _149_\[6\] _132_\[6\] VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__nand2_1
XFILLER_108_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11153_ net17 _05190_ _05192_ _158_\[15\] VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__a22o_1
XFILLER_1_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10104_ _04436_ _03984_ _04365_ _04318_ _04157_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__a311oi_2
X_11084_ net35 _01325_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__nor2_4
X_10035_ _142_\[21\] _04410_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11986_ _05982_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13725_ clknet_leaf_57_clk _00944_ VGND VGND VPWR VPWR _134_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10937_ net39 _04853_ _05098_ _05067_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__o211a_1
XFILLER_140_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13656_ clknet_leaf_56_clk _00875_ VGND VGND VPWR VPWR _138_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12607_ _06342_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__clkbuf_1
X_10868_ _05028_ _05049_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__or2_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13587_ clknet_leaf_46_clk _00806_ VGND VGND VPWR VPWR _142_\[19\] sky130_fd_sc_hd__dfxtp_1
X_10799_ _01418_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12538_ _06306_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12469_ _06270_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06961_ _01568_ _01570_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__or2_1
X_09680_ _185_\[6\] _03869_ _03919_ _04071_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__o211a_1
X_08700_ _01355_ _03118_ _03126_ _02355_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__a211o_1
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06892_ _179_\[31\] _01269_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__and2_1
X_08631_ _03056_ _03059_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08562_ _02990_ _02992_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07513_ _01684_ _02062_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__xnor2_1
X_08493_ _02878_ _02899_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__nor2_1
X_07444_ _182_\[10\] _01635_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__or2_1
XFILLER_90_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07375_ _185_\[8\] _234_\[8\] VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__or2_1
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09114_ _03516_ _03527_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09045_ _03426_ _03432_ _03459_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09947_ _04299_ _04306_ _142_\[16\] _04298_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09878_ _04252_ _04261_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__and2_1
XFILLER_85_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08829_ _03233_ _03235_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__nand2_1
XFILLER_45_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11840_ _05836_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__or2_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11771_ _05785_ _05786_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__and2_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13510_ clknet_leaf_60_clk _00729_ VGND VGND VPWR VPWR _152_\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _173_\[14\] _04917_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__or2_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10653_ _173_\[25\] _176_\[25\] _01226_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__mux2_1
X_13441_ clknet_leaf_122_clk _00660_ VGND VGND VPWR VPWR _164_\[27\] sky130_fd_sc_hd__dfxtp_1
X_10584_ _173_\[2\] _04849_ _04851_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__a21o_1
X_13372_ clknet_leaf_126_clk _00591_ VGND VGND VPWR VPWR _170_\[22\] sky130_fd_sc_hd__dfxtp_1
X_12323_ _06193_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12254_ _06157_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__clkbuf_1
X_11205_ _152_\[3\] _01368_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__and2_1
X_12185_ _140_\[20\] _138_\[20\] _06112_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__mux2_1
XFILLER_110_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11136_ _01259_ _05230_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__nand2_1
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11067_ _164_\[27\] _04872_ _04633_ _05181_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__o211a_1
X_10018_ _04345_ _04346_ _04372_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__and3_1
XFILLER_91_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11969_ _152_\[22\] _05965_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__or2_1
X_13708_ clknet_leaf_77_clk _00927_ VGND VGND VPWR VPWR _134_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13639_ clknet_leaf_53_clk _00858_ VGND VGND VPWR VPWR _138_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07160_ _237_\[0\] _01723_ _01411_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__mux2_1
X_07091_ _173_\[19\] _01667_ _01617_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__mux2_1
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09801_ _142_\[11\] _04187_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__and2_1
X_09732_ _04120_ _04121_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__or2_1
XFILLER_115_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07993_ _02527_ _02441_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__and2b_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06944_ _01420_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__clkbuf_4
X_09663_ _01241_ _01280_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__nor2_2
X_06875_ _243_\[27\] _01474_ _01461_ _01507_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__o211a_1
XFILLER_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09594_ _03973_ _03988_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08614_ _01847_ _03011_ _03042_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__a21oi_4
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _02940_ _02975_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__nand2_1
XFILLER_36_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_128_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_128_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08476_ _01710_ _02909_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__or2_1
X_07427_ _01978_ _01979_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__nand2_1
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07358_ _01856_ _01892_ _01914_ _01884_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__a211o_1
XFILLER_50_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07289_ _01846_ _01847_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09028_ _02839_ _03443_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__xnor2_2
XFILLER_104_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12941_ clknet_leaf_39_clk _00160_ VGND VGND VPWR VPWR _246_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12872_ _118_\[27\] _120_\[27\] _06473_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__mux2_1
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _140_\[19\] _05833_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_119_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_119_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _05769_ _05770_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__or2b_1
XFILLER_121_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _149_\[27\] _05709_ _05625_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__mux2_1
X_10705_ _167_\[9\] _04925_ _04933_ _04891_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__o211a_1
X_13424_ clknet_leaf_1_clk _00643_ VGND VGND VPWR VPWR _164_\[10\] sky130_fd_sc_hd__dfxtp_2
X_10636_ _173_\[20\] _176_\[20\] _01226_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__mux2_1
X_13355_ clknet_leaf_12_clk _00574_ VGND VGND VPWR VPWR _170_\[5\] sky130_fd_sc_hd__dfxtp_1
X_10567_ _176_\[29\] _179_\[29\] _04830_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__mux2_1
XFILLER_10_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10498_ _176_\[9\] _179_\[9\] _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__mux2_1
X_12306_ _06184_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__clkbuf_1
X_13286_ clknet_leaf_24_clk _00505_ VGND VGND VPWR VPWR _176_\[0\] sky130_fd_sc_hd__dfxtp_1
X_12237_ _06148_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12168_ _01393_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__clkbuf_4
X_12099_ _140_\[11\] _142_\[11\] _06068_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__mux2_1
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11119_ _158_\[7\] _01256_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 din[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_4
X_06660_ _01308_ _01340_ _01357_ _01303_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__o31a_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06591_ net35 VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08330_ _225_\[7\] VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_60_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08261_ _02686_ _02739_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__or2_1
XFILLER_20_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07212_ _182_\[3\] _01612_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__nand2_1
XFILLER_20_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08192_ _01406_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07143_ _173_\[31\] _01646_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__or2_1
XFILLER_145_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07074_ _173_\[15\] _01654_ _01617_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07976_ _02488_ _02489_ _02510_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__a21oi_1
X_09715_ _01281_ _03960_ _04080_ _04075_ _03872_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__a221oi_1
X_06927_ _176_\[9\] _240_\[9\] _01449_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__mux2_1
XFILLER_28_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09646_ _03998_ _04022_ _04037_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__o21bai_1
XFILLER_83_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06858_ _01495_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09577_ _185_\[2\] _03869_ _03919_ _03972_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__o211a_1
X_06789_ _01412_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08528_ _02957_ _02959_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__xnor2_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08459_ _185_\[1\] _02892_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11470_ _118_\[9\] _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10421_ _179_\[19\] _182_\[19\] _04693_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__mux2_1
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13140_ clknet_4_2_0_clk _00359_ VGND VGND VPWR VPWR _228_\[20\] sky130_fd_sc_hd__dfxtp_1
X_10352_ _04685_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13071_ clknet_leaf_107_clk _00290_ VGND VGND VPWR VPWR _234_\[15\] sky130_fd_sc_hd__dfxtp_1
X_12022_ net19 _06015_ _05785_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__mux2_1
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10283_ _179_\[5\] _04638_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__or2_1
XFILLER_2_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13973_ clknet_leaf_93_clk _01192_ VGND VGND VPWR VPWR _118_\[21\] sky130_fd_sc_hd__dfxtp_2
XFILLER_19_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12924_ clknet_leaf_28_clk _436_\[1\] _00101_ VGND VGND VPWR VPWR _392_\[1\] sky130_fd_sc_hd__dfstp_2
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _118_\[19\] _120_\[19\] _06462_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__mux2_1
XFILLER_34_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11806_ _05804_ _05808_ _05817_ _05776_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__a31oi_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12786_ _06436_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__clkbuf_1
X_11737_ _05755_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__clkbuf_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11668_ _116_\[26\] _05693_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__nand2_1
XFILLER_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10619_ _02085_ _04861_ _04875_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__a21boi_1
X_11599_ _05612_ _05614_ _05622_ _05632_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__o31a_1
X_13407_ clknet_leaf_127_clk _00626_ VGND VGND VPWR VPWR _167_\[25\] sky130_fd_sc_hd__dfxtp_2
X_13338_ clknet_leaf_0_clk _00557_ VGND VGND VPWR VPWR _173_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13269_ clknet_leaf_25_clk _00488_ VGND VGND VPWR VPWR _179_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07830_ _02368_ _02369_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__or2_1
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07761_ _01694_ _02302_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__xnor2_2
X_09500_ _01280_ _03897_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__nand2_2
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06712_ _01388_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07692_ _02227_ _02229_ _02226_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__a21oi_2
X_06643_ _01306_ _01344_ _01268_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__o21a_1
XFILLER_92_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09431_ _03834_ _03835_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__xor2_1
X_06574_ _01282_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__clkbuf_4
X_09362_ _170_\[27\] _02858_ _03702_ _03767_ _03768_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__a221o_1
XFILLER_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08313_ _02776_ _02733_ _02760_ _02777_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__o211a_1
XANTENNA_11 _128_\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _179_\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09293_ _03599_ _03663_ _03664_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__a21boi_1
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_33 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08244_ _231_\[15\] _02690_ _02712_ _02727_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__a211o_1
XANTENNA_44 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _173_\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08175_ _02625_ _02677_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__or2_1
XFILLER_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_88 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07126_ _01420_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07057_ _240_\[11\] _01583_ _01607_ _01641_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__a211o_1
XFILLER_133_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07959_ _243_\[27\] _240_\[27\] _01694_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__mux2_4
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10970_ _01435_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__buf_4
XFILLER_16_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09629_ _04000_ _04014_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__nor2_1
XFILLER_43_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12640_ _126_\[12\] _124_\[12\] _06357_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__mux2_1
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_16
X_12571_ _06323_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11522_ _149_\[10\] _05563_ _05533_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__mux2_1
XFILLER_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11453_ _05496_ _05498_ _05495_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__a21oi_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10404_ _176_\[14\] _04683_ _04723_ _01419_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__a211o_1
X_11384_ _05435_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__inv_2
X_13123_ clknet_leaf_116_clk _00342_ VGND VGND VPWR VPWR _228_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10335_ _182_\[27\] _04654_ _04671_ _01710_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__a31o_1
XFILLER_133_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10266_ _182_\[0\] _01218_ _04631_ _03309_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__a31o_1
XFILLER_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13054_ clknet_leaf_110_clk _00273_ VGND VGND VPWR VPWR _237_\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12005_ _05986_ _05991_ _05984_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__o21ai_1
XFILLER_105_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10197_ _04565_ _04566_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13956_ clknet_leaf_71_clk _01175_ VGND VGND VPWR VPWR _118_\[4\] sky130_fd_sc_hd__dfxtp_2
X_13887_ clknet_leaf_69_clk _01106_ VGND VGND VPWR VPWR _124_\[31\] sky130_fd_sc_hd__dfxtp_1
X_12907_ clknet_leaf_86_clk _00131_ VGND VGND VPWR VPWR _116_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12838_ _06463_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__clkbuf_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12769_ _06427_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_41_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput31 din[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 din[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09980_ _04082_ _04320_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__nor2_1
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08931_ _03347_ _03348_ _02161_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08862_ _02064_ _03255_ _03282_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__o21a_1
XFILLER_84_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07813_ _01437_ _02353_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__and2_1
XFILLER_123_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08793_ _03208_ _03209_ _03216_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__o21ai_1
X_07744_ _02172_ _02286_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__or2_1
XFILLER_37_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07675_ _02218_ _02219_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__and2_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06626_ _392_\[1\] _392_\[0\] _01210_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__a21oi_1
X_09414_ _03817_ _03818_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__nand2_1
XFILLER_25_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06557_ _158_\[21\] _01265_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_32_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
X_09345_ _03750_ _03751_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__and2_1
X_09276_ _03683_ _03684_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__or2_1
XFILLER_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08227_ _02686_ _02715_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__or2_1
XFILLER_107_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08158_ _234_\[22\] _02646_ _02664_ _02666_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__a211o_1
XFILLER_134_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07109_ _173_\[23\] _01681_ _01672_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__mux2_1
X_08089_ _167_\[3\] _02616_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__or2_1
X_10120_ _03946_ _04492_ _04493_ _00105_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__o211a_1
XFILLER_106_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10051_ _04395_ _04405_ _04393_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__o21ba_1
XFILLER_88_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13810_ clknet_leaf_94_clk _01029_ VGND VGND VPWR VPWR _128_\[18\] sky130_fd_sc_hd__dfxtp_1
X_13741_ clknet_leaf_80_clk _00960_ VGND VGND VPWR VPWR _132_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10953_ net44 _05068_ _05109_ _05086_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__a211o_1
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13672_ clknet_leaf_54_clk _00891_ VGND VGND VPWR VPWR _136_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10884_ _167_\[29\] _05059_ _05043_ _05060_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__o211a_1
X_12623_ _126_\[4\] _124_\[4\] _06346_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_23_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_71_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12554_ _128_\[3\] _126_\[3\] _06313_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__mux2_1
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11505_ _118_\[12\] _05547_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12485_ _06278_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11436_ _116_\[2\] _05485_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__and2_1
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11367_ _149_\[25\] _132_\[25\] VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__nand2_1
XFILLER_98_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10318_ _179_\[19\] _04646_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__or2_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13106_ clknet_leaf_117_clk _00325_ VGND VGND VPWR VPWR _231_\[18\] sky130_fd_sc_hd__dfxtp_1
X_11298_ _152_\[15\] _05366_ _05318_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__mux2_1
X_13037_ clknet_leaf_81_clk _00256_ VGND VGND VPWR VPWR _237_\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ _01244_ _01285_ _03952_ _01239_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__a211o_1
XFILLER_78_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13939_ clknet_leaf_96_clk _01158_ VGND VGND VPWR VPWR _120_\[19\] sky130_fd_sc_hd__dfxtp_1
X_07460_ _02010_ _02011_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__nand2_1
X_07391_ _01520_ _01922_ _01945_ _01946_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
X_09130_ _03476_ _03542_ _03509_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__o21a_1
X_09061_ _03469_ _03475_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__and2b_1
XFILLER_135_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08012_ _02544_ _02545_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__nor2_1
XFILLER_143_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09963_ _04326_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__inv_2
XFILLER_103_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08914_ _170_\[15\] _02817_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__nor2_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09894_ _04275_ _04276_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__or2_1
XFILLER_97_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08845_ _03252_ _03266_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__xor2_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08776_ _01985_ _03163_ _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__a21oi_2
XFILLER_57_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07727_ _02268_ _02269_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__or2_1
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07658_ _01661_ _01827_ _02178_ _02203_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__a211o_1
XFILLER_13_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06609_ _01246_ _01268_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__nor2_1
X_07589_ _02135_ _02136_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__and2b_1
XFILLER_40_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_clk clknet_3_4_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09328_ _02404_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__nand2_1
XFILLER_138_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09259_ _02380_ _03662_ _03668_ _01439_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__o211a_1
X_12270_ _06165_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11221_ _149_\[6\] _132_\[6\] VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__or2_1
XFILLER_135_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11152_ _01262_ _05242_ _05194_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10103_ _03886_ _03976_ _04476_ _01233_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__o31a_1
XFILLER_1_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11083_ _03866_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__inv_2
X_10034_ _142_\[21\] _04410_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__and2_1
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11985_ _142_\[23\] _05981_ _05893_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__mux2_1
XFILLER_56_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13724_ clknet_leaf_57_clk _00943_ VGND VGND VPWR VPWR _134_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10936_ _05079_ _05097_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__or2_1
X_13655_ clknet_leaf_48_clk _00874_ VGND VGND VPWR VPWR _138_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10867_ _167_\[24\] _170_\[24\] _04995_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__mux2_1
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _128_\[28\] _126_\[28\] _06335_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__mux2_1
XFILLER_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13586_ clknet_leaf_46_clk _00805_ VGND VGND VPWR VPWR _142_\[18\] sky130_fd_sc_hd__dfxtp_1
X_10798_ _167_\[4\] _04980_ _04958_ _04999_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__o211a_1
XFILLER_118_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12537_ _130_\[27\] _128_\[27\] _06302_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__mux2_1
XFILLER_8_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12468_ _132_\[26\] _130_\[26\] _06269_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__mux2_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11419_ _149_\[31\] _132_\[31\] VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12399_ _132_\[25\] _134_\[25\] _06230_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__mux2_1
XFILLER_113_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06960_ _176_\[18\] _240_\[18\] _01569_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_3_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_39_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06891_ _01519_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__buf_4
XFILLER_67_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08630_ _03025_ _03058_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__nand2_1
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08561_ _228_\[4\] _231_\[4\] _02991_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__o21a_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07512_ _01667_ _01623_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__xnor2_1
X_08492_ _02922_ _02924_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__xnor2_2
X_07443_ _182_\[10\] _01635_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__nand2_1
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07374_ _01667_ _01929_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__xnor2_2
XFILLER_50_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09113_ _02311_ _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09044_ _03426_ _03432_ _03459_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__and3_1
XFILLER_135_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09946_ _04324_ _04326_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09877_ _04161_ _04254_ _04260_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__o21ai_1
XFILLER_97_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08828_ _02807_ _02845_ _02834_ _03250_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__o211a_1
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08759_ _03181_ _03183_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__xor2_2
X_11770_ _05777_ _05783_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__nand2_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10721_ _04682_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__buf_2
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ clknet_leaf_127_clk _00659_ VGND VGND VPWR VPWR _164_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10652_ _04855_ _04896_ _04897_ _04839_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__a211o_1
XFILLER_9_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10583_ _176_\[2\] net68 _01751_ _04682_ _02711_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__a221o_1
X_13371_ clknet_leaf_130_clk _00590_ VGND VGND VPWR VPWR _170_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12322_ _136_\[21\] _134_\[21\] _06189_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__mux2_1
XFILLER_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12253_ _138_\[20\] _136_\[20\] _06156_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__mux2_1
X_11204_ _05274_ _05283_ _05282_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__o21ai_1
XFILLER_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12184_ _06120_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11135_ _158_\[10\] _01258_ _158_\[11\] VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11066_ _03735_ _04681_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10017_ _04393_ _04394_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__or2b_1
XFILLER_76_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13707_ clknet_leaf_48_clk _00926_ VGND VGND VPWR VPWR _134_\[11\] sky130_fd_sc_hd__dfxtp_1
X_11968_ _152_\[22\] _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__nand2_1
XFILLER_60_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11899_ _140_\[26\] _05902_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__xnor2_2
X_10919_ _01418_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__buf_2
X_13638_ clknet_leaf_53_clk _00857_ VGND VGND VPWR VPWR _138_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13569_ clknet_leaf_54_clk _00788_ VGND VGND VPWR VPWR _142_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07090_ _237_\[19\] VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__buf_6
XFILLER_8_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09800_ _246_\[11\] _01314_ _03914_ _243_\[11\] _01464_ VGND VGND VPWR VPWR _04187_
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07992_ _02474_ _02473_ _02481_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__or3_1
X_09731_ _04119_ _04101_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__and2b_1
XFILLER_101_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06943_ _01435_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__clkbuf_4
XFILLER_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09662_ _01230_ _03933_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__nor2_1
X_06874_ _179_\[27\] _01301_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__or2_1
XFILLER_95_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09593_ _03975_ _03987_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__xor2_1
XFILLER_131_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08613_ _03008_ _03010_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__nor2_1
XFILLER_67_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _02932_ _02934_ _02941_ _02943_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__o211ai_1
XFILLER_63_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08475_ _02772_ _02908_ _01411_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__mux2_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07426_ _185_\[10\] _234_\[10\] VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__nand2_1
XFILLER_50_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07357_ _01911_ _01912_ _01913_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07288_ _243_\[5\] _240_\[5\] _01620_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__mux2_4
X_09027_ _02797_ _02768_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09929_ _04295_ _04296_ _04310_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__a21o_1
XFILLER_58_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12940_ clknet_leaf_40_clk _00159_ VGND VGND VPWR VPWR _246_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12871_ _06480_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _140_\[26\] _140_\[28\] VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _152_\[3\] _05768_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__or2_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11684_ _05707_ _05708_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__xnor2_1
X_10704_ _04888_ _04932_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__or2_1
XFILLER_139_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10635_ _173_\[19\] _04848_ _04885_ _04839_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__a211o_1
X_13423_ clknet_leaf_2_clk _00642_ VGND VGND VPWR VPWR _164_\[9\] sky130_fd_sc_hd__dfxtp_1
X_13354_ clknet_leaf_11_clk _00573_ VGND VGND VPWR VPWR _170_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12305_ _136_\[13\] _134_\[13\] _06178_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__mux2_1
X_10566_ _173_\[28\] _04836_ _04838_ _04839_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__a211o_1
XFILLER_127_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13285_ clknet_leaf_5_clk _00504_ VGND VGND VPWR VPWR _179_\[31\] sky130_fd_sc_hd__dfxtp_1
X_10497_ _01214_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__buf_4
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12236_ _138_\[12\] _136_\[12\] _06145_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__mux2_1
X_12167_ _06111_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11118_ _05217_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12098_ _06075_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11049_ _164_\[20\] _01218_ _04648_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__o21a_1
Xinput7 din[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XFILLER_92_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06590_ _01276_ _01292_ _01294_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__a21oi_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08260_ _164_\[20\] _228_\[20\] _02687_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__mux2_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07211_ _182_\[3\] _01612_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__nor2_1
X_08191_ _231_\[0\] _02659_ _02636_ _02689_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__o211a_1
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07142_ _237_\[31\] VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__buf_6
XFILLER_20_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07073_ _237_\[15\] VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__clkbuf_4
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07975_ _02506_ _02509_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__xor2_1
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09714_ _04103_ _04080_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__or2_1
X_06926_ _01480_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__buf_2
XFILLER_28_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09645_ _03998_ _04022_ _04037_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__or3b_1
X_06857_ _01405_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__buf_4
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09576_ _03970_ _03971_ _03946_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__a21o_1
X_06788_ _246_\[4\] _01407_ _01436_ _01443_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__a211o_1
XFILLER_82_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08527_ _01762_ _02918_ _02958_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__a21oi_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08458_ _02846_ _02891_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__xnor2_2
X_07409_ _01936_ _01950_ _01961_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10420_ _04671_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08389_ net48 _02835_ _01353_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__mux2_1
XFILLER_136_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10351_ _04625_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__buf_2
X_10282_ _179_\[4\] _04629_ _04643_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__a21o_1
X_13070_ clknet_leaf_83_clk _00289_ VGND VGND VPWR VPWR _234_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12021_ _06010_ _06014_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__xor2_1
XFILLER_105_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13972_ clknet_leaf_93_clk _01191_ VGND VGND VPWR VPWR _118_\[20\] sky130_fd_sc_hd__dfxtp_2
X_12923_ clknet_leaf_32_clk _436_\[0\] _00100_ VGND VGND VPWR VPWR _392_\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_19_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12854_ _06471_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11805_ _05804_ _05808_ _05817_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__a21o_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12785_ _122_\[17\] _120_\[17\] _06434_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__mux2_1
X_11736_ _142_\[1\] _05754_ _05625_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__mux2_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11667_ _118_\[12\] _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10618_ _176_\[13\] _04678_ _04627_ _173_\[13\] _02833_ VGND VGND VPWR VPWR _04875_
+ sky130_fd_sc_hd__o221a_1
X_11598_ _05610_ _05619_ _05620_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__a21o_1
X_13406_ clknet_leaf_126_clk _00625_ VGND VGND VPWR VPWR _167_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10549_ _176_\[24\] _04771_ _04806_ _04826_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__o211a_1
X_13337_ clknet_leaf_10_clk _00556_ VGND VGND VPWR VPWR _173_\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13268_ clknet_leaf_24_clk _00487_ VGND VGND VPWR VPWR _179_\[14\] sky130_fd_sc_hd__dfxtp_1
X_12219_ _138_\[4\] _136_\[4\] _06134_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__mux2_1
X_13199_ clknet_leaf_34_clk _00418_ VGND VGND VPWR VPWR _185_\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_123_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_07760_ _01650_ _237_\[0\] VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__xnor2_2
XFILLER_56_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06711_ _118_\[20\] _116_\[20\] _01381_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__mux2_1
XFILLER_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07691_ _02233_ _02234_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__and2b_2
X_09430_ _03762_ _03765_ _03800_ _03802_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__a31o_1
XFILLER_25_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06642_ _096_ _01208_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__nand2_1
XFILLER_80_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06573_ _195_\[0\] VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__clkbuf_4
X_09361_ _170_\[27\] _02858_ _02855_ _170_\[26\] VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__o211a_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09292_ _03600_ _03606_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__nor2_1
XFILLER_21_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08312_ net58 _02736_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__or2_1
XFILLER_33_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_12 _142_\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_23 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08243_ _228_\[15\] _02698_ _02723_ _02726_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__o211a_1
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_34 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_78 _179_\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08174_ _167_\[28\] _231_\[28\] _02626_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__mux2_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_89 _173_\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07125_ _237_\[27\] VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__buf_4
XFILLER_134_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07056_ _01638_ _01639_ _01609_ _01640_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__o211a_1
XFILLER_133_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07958_ _02492_ _02493_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__or2_1
X_06909_ _243_\[3\] _01496_ _01509_ _01533_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__a211o_1
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07889_ _02425_ _02426_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__nand2_1
X_09628_ _185_\[4\] _03869_ _03919_ _04021_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__o211a_1
XFILLER_55_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09559_ _03954_ _03901_ _03938_ _03935_ _03879_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__a32o_1
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12570_ _128_\[11\] _126_\[11\] _06313_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__mux2_1
XFILLER_141_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11521_ _05560_ _05562_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__xor2_1
XFILLER_11_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11452_ _05500_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11383_ _05440_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__clkbuf_1
X_10403_ _179_\[14\] _04721_ _04705_ _04722_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__o211a_1
X_10334_ _182_\[26\] _04663_ _04673_ _04649_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__o211a_1
X_13122_ clknet_leaf_115_clk _00341_ VGND VGND VPWR VPWR _228_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13053_ clknet_leaf_108_clk _00272_ VGND VGND VPWR VPWR _237_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__buf_4
X_10196_ _142_\[27\] _04538_ _04539_ _04546_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__o2bb2a_1
X_12004_ _05997_ _05998_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__or2_1
XFILLER_87_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13955_ clknet_leaf_71_clk _01174_ VGND VGND VPWR VPWR _118_\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_81_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13886_ clknet_leaf_69_clk _01105_ VGND VGND VPWR VPWR _124_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12906_ clknet_leaf_86_clk _00130_ VGND VGND VPWR VPWR _116_\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _118_\[10\] _120_\[10\] _06462_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__mux2_1
XFILLER_34_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12768_ _122_\[9\] _120_\[9\] _06423_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__mux2_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12699_ _124_\[8\] _122_\[8\] _06390_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__mux2_1
X_11719_ _05737_ _05739_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput10 din[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 din[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
XFILLER_30_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput32 din[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08930_ _02161_ _03347_ _03348_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__and3_1
XFILLER_123_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08861_ _185_\[13\] _03254_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__nand2_1
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07812_ _02350_ _02352_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__xor2_2
X_08792_ _01778_ _03215_ _01412_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__o21a_1
XFILLER_38_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07743_ _02170_ _02179_ _02227_ _02235_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__or4bb_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07674_ _02189_ _02204_ _02217_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__or3_1
XFILLER_25_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06625_ _01207_ _01208_ _01268_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__nor3_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09413_ _185_\[30\] _03816_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__or2_1
XFILLER_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06556_ _158_\[19\] _158_\[20\] _01264_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__or3_1
X_09344_ _03714_ _03743_ _03749_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__nand3_1
XFILLER_21_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09275_ _03647_ _03671_ _03682_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__and3_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08226_ _164_\[10\] _228_\[10\] _02687_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__mux2_1
X_08157_ _231_\[22\] _02649_ _02641_ _02665_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__o211a_1
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07108_ _237_\[23\] VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__buf_6
X_08088_ _01339_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__clkbuf_2
XFILLER_121_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07039_ _01626_ _01565_ _01609_ _01627_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__o211a_1
X_10050_ _04425_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__and2b_1
XFILLER_0_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13740_ clknet_leaf_78_clk _00959_ VGND VGND VPWR VPWR _132_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10952_ _164_\[17\] _05107_ _05094_ _05108_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__o211a_1
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13671_ clknet_leaf_54_clk _00890_ VGND VGND VPWR VPWR _136_\[7\] sky130_fd_sc_hd__dfxtp_1
X_10883_ _170_\[29\] _05036_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__or2_1
X_12622_ _06350_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12553_ _06314_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11504_ _118_\[27\] _118_\[16\] VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__xnor2_1
X_12484_ _130_\[2\] _128_\[2\] _06269_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__mux2_1
X_11435_ _118_\[20\] _05484_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11366_ _05425_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11297_ _05362_ _05365_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__xnor2_1
X_10317_ _182_\[18\] _04663_ _04664_ _04649_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__o211a_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13105_ clknet_leaf_117_clk _00324_ VGND VGND VPWR VPWR _231_\[17\] sky130_fd_sc_hd__dfxtp_1
X_10248_ _04132_ _04437_ _03950_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__or3b_1
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13036_ clknet_opt_1_0_clk _00255_ VGND VGND VPWR VPWR _237_\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10179_ _04548_ _04549_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__nor2_1
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13938_ clknet_leaf_96_clk _01157_ VGND VGND VPWR VPWR _120_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13869_ clknet_leaf_97_clk _01088_ VGND VGND VPWR VPWR _124_\[13\] sky130_fd_sc_hd__dfxtp_1
X_07390_ _01943_ _01924_ _01925_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__or3_1
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09060_ _03375_ _03470_ _03474_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__o21ai_1
XFILLER_135_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08011_ _02506_ _02508_ _02507_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__a21boi_1
XFILLER_128_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09962_ _04339_ _04341_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__xor2_1
XFILLER_104_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08913_ _03310_ _03311_ _03331_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__a21oi_1
XFILLER_131_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09893_ _142_\[15\] _04274_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__nor2_1
XFILLER_69_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08844_ _03263_ _03265_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__xnor2_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ _03160_ _03162_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__nor2_1
XFILLER_73_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07726_ _02244_ _02246_ _02267_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__and3_1
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07657_ _01520_ _02181_ _02201_ _02202_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__o211a_1
X_06608_ _01208_ _01250_ _01310_ _01295_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__o211a_1
X_07588_ _182_\[15\] _01654_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__nand2_1
XFILLER_43_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06539_ _01206_ _01247_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__or2_2
X_09327_ _03733_ _03734_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__xor2_2
XFILLER_139_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09258_ _01519_ _03667_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__or2_1
XFILLER_135_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08209_ _228_\[5\] _02698_ _02679_ _02702_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__o211a_1
X_09189_ _03598_ _03599_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__nand2_1
XFILLER_4_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11220_ _05298_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11151_ _158_\[15\] _01261_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__nand2_1
XFILLER_134_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10102_ _01292_ _04057_ _04475_ _01238_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11082_ _03866_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__inv_2
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10033_ _246_\[21\] _01315_ _04409_ _243_\[21\] _01493_ VGND VGND VPWR VPWR _04410_
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11984_ net16 _05980_ _05785_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__mux2_1
X_13723_ clknet_leaf_57_clk _00942_ VGND VGND VPWR VPWR _134_\[27\] sky130_fd_sc_hd__dfxtp_1
X_10935_ _164_\[12\] _167_\[12\] _05064_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__mux2_1
X_13654_ clknet_leaf_56_clk _00873_ VGND VGND VPWR VPWR _138_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10866_ _04671_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__buf_4
XFILLER_32_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12605_ _06341_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__clkbuf_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13585_ clknet_leaf_45_clk _00804_ VGND VGND VPWR VPWR _142_\[17\] sky130_fd_sc_hd__dfxtp_1
X_10797_ _170_\[4\] _04953_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__or2_1
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12536_ _06305_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12467_ _06200_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__clkbuf_4
XFILLER_138_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11418_ _05465_ _05468_ _05464_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__a21o_1
XFILLER_125_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12398_ _06233_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11349_ _05410_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__inv_2
XFILLER_4_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06890_ _01518_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__buf_4
X_13019_ clknet_leaf_13_clk _00238_ VGND VGND VPWR VPWR _240_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08560_ _228_\[4\] _231_\[4\] _02781_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__a21o_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07511_ _02047_ _02048_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__and2b_1
X_08491_ _228_\[2\] _231_\[2\] _02923_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__o21a_1
X_07442_ _01991_ _01993_ _01409_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__a21oi_1
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07373_ _01650_ _01604_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09112_ _03519_ _03525_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__xor2_1
XFILLER_129_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09043_ _03457_ _03458_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__and2b_1
XFILLER_129_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09945_ _142_\[17\] _04325_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09876_ _04255_ _04256_ _04257_ _04259_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__o211a_1
XFILLER_58_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08827_ _01355_ _03241_ _03242_ _03249_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__a31o_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08758_ _03129_ _03131_ _03182_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__a21oi_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08689_ _03081_ _03082_ _03083_ _03080_ _03078_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__o32a_1
X_07709_ _02251_ _02252_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10720_ _167_\[13\] _04836_ _04944_ _04914_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__a211o_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10651_ _02416_ _04631_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__nor2_1
X_10582_ _173_\[1\] _04849_ _04850_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__a21o_1
XFILLER_70_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13370_ clknet_leaf_130_clk _00589_ VGND VGND VPWR VPWR _170_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12321_ _06192_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12252_ _01393_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__clkbuf_4
XFILLER_135_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11203_ _05274_ _05282_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__or3_1
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12183_ _140_\[19\] _138_\[19\] _06112_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__mux2_1
X_11134_ _05227_ _05228_ _05229_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__a21o_1
XFILLER_96_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11065_ _03704_ _04855_ _04628_ net54 _05180_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__o221a_1
XFILLER_1_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10016_ _04356_ _04376_ _04392_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__or3b_1
XFILLER_95_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11967_ _140_\[7\] _140_\[9\] VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__xor2_2
XFILLER_51_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13706_ clknet_leaf_48_clk _00925_ VGND VGND VPWR VPWR _134_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10918_ _164_\[7\] _05059_ _05043_ _05084_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__o211a_1
X_11898_ _140_\[1\] _140_\[3\] VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__xnor2_2
X_13637_ clknet_leaf_54_clk _00856_ VGND VGND VPWR VPWR _138_\[5\] sky130_fd_sc_hd__dfxtp_1
X_10849_ _01216_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__clkbuf_2
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13568_ clknet_leaf_55_clk _00787_ VGND VGND VPWR VPWR _142_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12519_ _06296_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13499_ clknet_leaf_36_clk _00718_ VGND VGND VPWR VPWR _158_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07991_ _02524_ _02525_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__nor2_1
X_09730_ _04101_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__and2b_1
Xclkbuf_4_7_0_clk clknet_3_3_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_06942_ _243_\[13\] _01548_ _01545_ _01556_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__o211a_1
XFILLER_86_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09661_ _04028_ _04050_ _04052_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__a21bo_1
X_06873_ _246_\[26\] _01485_ _01481_ _01506_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__o211a_1
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09592_ _03978_ _03980_ _03986_ _03910_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__a2bb2o_1
X_08612_ _01875_ _03040_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__xnor2_4
XFILLER_54_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08543_ _02972_ _02973_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__and2b_1
XFILLER_63_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08474_ _02904_ _02905_ _01269_ _02907_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07425_ _185_\[10\] _234_\[10\] VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__or2_1
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07356_ _01911_ _01912_ _01523_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__o21ai_1
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07287_ _01844_ _01845_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__or2_1
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09026_ _03422_ _03424_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__and2b_1
XFILLER_123_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09928_ _04308_ _04309_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__nand2_1
XFILLER_49_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09859_ _04207_ _04219_ _04242_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__or3b_1
XFILLER_105_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _118_\[26\] _120_\[26\] _06473_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__mux2_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _142_\[8\] _05279_ _05832_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__o21a_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _152_\[3\] _05768_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__and2_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11683_ _05695_ _05700_ _05694_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__a21bo_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10703_ _170_\[9\] _173_\[9\] _04830_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__mux2_1
X_10634_ _176_\[19\] _04872_ _04633_ _04884_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__o211a_1
X_13422_ clknet_leaf_12_clk _00641_ VGND VGND VPWR VPWR _164_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13353_ clknet_leaf_2_clk _00572_ VGND VGND VPWR VPWR _170_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12304_ _06183_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__clkbuf_1
X_10565_ _01418_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__clkbuf_4
X_10496_ _173_\[8\] _04780_ _04789_ _04785_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__o211a_1
X_13284_ clknet_leaf_5_clk _00503_ VGND VGND VPWR VPWR _179_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12235_ _06147_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12166_ _140_\[11\] _138_\[11\] _06101_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__mux2_1
X_11117_ _05216_ _158_\[6\] _05192_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__mux2_1
XFILLER_96_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12097_ _140_\[10\] _142_\[10\] _06068_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__mux2_1
XFILLER_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11048_ net46 _04848_ _05170_ _01436_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__a211o_1
Xinput8 din[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_92_787 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12999_ clknet_leaf_15_clk _00218_ VGND VGND VPWR VPWR _240_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07210_ _01771_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08190_ _02686_ _02688_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__or2_1
X_07141_ _240_\[30\] _01660_ _01653_ _01706_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__o211a_1
XFILLER_145_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07072_ _01480_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07974_ _02507_ _02508_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__nand2_1
X_09713_ _04002_ _03901_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__nand2_2
X_06925_ _243_\[8\] _01536_ _01509_ _01544_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__a211o_1
X_09644_ _04035_ _04036_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__nand2_1
X_06856_ _246_\[21\] _01407_ _01460_ _01494_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__a211o_1
XFILLER_82_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09575_ _03968_ _03969_ _03943_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__o21ai_1
X_06787_ _243_\[4\] _01438_ _01439_ _01442_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__o211a_1
XFILLER_82_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08526_ _02915_ _02917_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__nor2_1
XFILLER_24_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08457_ _02814_ _225_\[3\] VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__xnor2_1
X_07408_ _01936_ _01950_ _01961_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__or3_1
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08388_ _225_\[20\] VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__clkbuf_4
XFILLER_137_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07339_ _01664_ _01895_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10350_ _01225_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__clkbuf_4
X_10281_ _182_\[4\] _01218_ _04642_ _03309_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__a31o_1
X_09009_ _03410_ _03411_ _03425_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__o21ai_1
XFILLER_117_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12020_ _05991_ _06011_ _06013_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__o21a_1
XFILLER_132_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13971_ clknet_leaf_96_clk _01190_ VGND VGND VPWR VPWR _118_\[19\] sky130_fd_sc_hd__dfxtp_2
X_12922_ clknet_leaf_88_clk _00146_ VGND VGND VPWR VPWR _116_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12853_ _118_\[18\] _120_\[18\] _06462_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__mux2_1
X_11804_ _05814_ _05816_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__nand2_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12784_ _06435_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ net12 _05753_ _05742_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__mux2_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11666_ _118_\[29\] _118_\[1\] VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__xnor2_1
X_13405_ clknet_leaf_128_clk _00624_ VGND VGND VPWR VPWR _167_\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10617_ _173_\[12\] _04849_ _04874_ _04839_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__a211o_1
X_11597_ _05629_ _05630_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__nand2_1
X_13336_ clknet_leaf_9_clk _00555_ VGND VGND VPWR VPWR _173_\[18\] sky130_fd_sc_hd__dfxtp_1
X_10548_ _179_\[24\] _04799_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__or2_1
XFILLER_6_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13267_ clknet_leaf_26_clk _00486_ VGND VGND VPWR VPWR _179_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12218_ _06138_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10479_ _173_\[3\] _04774_ _04776_ _04777_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__a211o_1
X_13198_ clknet_leaf_34_clk _00417_ VGND VGND VPWR VPWR _185_\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_123_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12149_ _06102_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06710_ _01387_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07690_ _182_\[19\] _01667_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__nand2_1
X_06641_ _01295_ _01342_ _01312_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__a21o_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06572_ _01280_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__clkbuf_4
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09360_ _03700_ _03733_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__nor2_1
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09291_ _03698_ _03699_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__nand2_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08311_ _225_\[2\] VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__buf_4
XFILLER_21_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08242_ _164_\[15\] _02701_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__or2_1
XANTENNA_13 _164_\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 _182_\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08173_ _234_\[27\] _02659_ _02636_ _02676_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__o211a_1
X_07124_ _01435_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__clkbuf_4
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07055_ _173_\[11\] _01580_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__or2_1
XFILLER_102_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07957_ _02453_ _02454_ _02491_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__and3_1
XFILLER_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06908_ _240_\[3\] _01526_ _01510_ _01532_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__o211a_1
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07888_ _02423_ _02424_ _02422_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__a21o_1
X_09627_ _04019_ _04020_ _03946_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__a21o_1
X_06839_ _179_\[17\] _01300_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__or2_1
XFILLER_71_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09558_ _01280_ _01282_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__nand2_1
XFILLER_12_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08509_ _170_\[3\] _225_\[3\] VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__nand2_1
X_09489_ _03884_ _03886_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__nor2_1
X_11520_ _05539_ _05544_ _05552_ _05561_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__o31a_1
XFILLER_51_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11451_ _149_\[3\] _05499_ _05439_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__mux2_1
XFILLER_109_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11382_ _152_\[26\] _05438_ _05439_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__mux2_1
X_10402_ _182_\[14\] _04696_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__or2_1
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10333_ _179_\[26\] _04646_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__or2_1
X_13121_ clknet_leaf_112_clk _00340_ VGND VGND VPWR VPWR _228_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13052_ clknet_leaf_110_clk _00271_ VGND VGND VPWR VPWR _237_\[28\] sky130_fd_sc_hd__dfxtp_1
X_10264_ _04625_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__buf_4
X_10195_ _04560_ _04564_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__xnor2_1
X_12003_ _05995_ _05996_ _152_\[25\] VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13954_ clknet_leaf_71_clk _01173_ VGND VGND VPWR VPWR _118_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13885_ clknet_leaf_72_clk _01104_ VGND VGND VPWR VPWR _124_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12905_ clknet_leaf_93_clk _00129_ VGND VGND VPWR VPWR _116_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12836_ _06004_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__buf_4
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12767_ _06426_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__clkbuf_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12698_ _01392_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__buf_6
X_11718_ _118_\[6\] _05738_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__xnor2_1
Xinput11 din[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 din[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
X_11649_ _118_\[10\] _05676_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__xnor2_1
Xinput33 dst_ready VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13319_ clknet_leaf_18_clk _00538_ VGND VGND VPWR VPWR _173_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08860_ _02124_ _03280_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07811_ _02291_ _02351_ _02297_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__o21a_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08791_ _03212_ _03214_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__xnor2_2
X_07742_ _02283_ _02233_ _02234_ _02284_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__o211a_1
XFILLER_38_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07673_ _02189_ _02204_ _02217_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__o21ai_1
X_06624_ _01246_ _01306_ _01316_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09412_ _185_\[30\] _03816_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__nand2_1
XFILLER_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09343_ _03714_ _03743_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__a21o_1
X_06555_ _158_\[18\] _01263_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__or2_1
XFILLER_33_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09274_ _03647_ _03671_ _03682_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08225_ _231_\[9\] _02690_ _02712_ _02714_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__a211o_1
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08156_ _167_\[22\] _02652_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__or2_1
XFILLER_5_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07107_ _240_\[22\] _01660_ _01653_ _01680_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__o211a_1
X_08087_ _234_\[2\] _02448_ _02419_ _02615_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__o211a_1
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07038_ _173_\[7\] _01580_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__or2_1
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08989_ _03405_ _03406_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__xor2_2
XFILLER_91_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10951_ _167_\[17\] _05089_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__or2_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13670_ clknet_leaf_54_clk _00889_ VGND VGND VPWR VPWR _136_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12621_ _126_\[3\] _124_\[3\] _06346_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__mux2_1
XFILLER_73_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10882_ _01225_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__clkbuf_4
XFILLER_52_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12552_ _128_\[2\] _126_\[2\] _06313_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__mux2_1
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12483_ _06277_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__clkbuf_1
X_11503_ _05546_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11434_ _118_\[9\] _118_\[5\] VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11365_ _152_\[24\] _05424_ _05318_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_100_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_100_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11296_ _05355_ _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__nand2_1
X_10316_ _179_\[18\] _04646_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__or2_1
X_13104_ clknet_leaf_105_clk _00323_ VGND VGND VPWR VPWR _231_\[16\] sky130_fd_sc_hd__dfxtp_1
X_10247_ _04055_ _04077_ _04361_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__or3_1
X_13035_ clknet_leaf_45_clk _00254_ VGND VGND VPWR VPWR _237_\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10178_ _04515_ _04524_ _04547_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__o21ba_1
XFILLER_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13937_ clknet_leaf_95_clk _01156_ VGND VGND VPWR VPWR _120_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13868_ clknet_leaf_97_clk _01087_ VGND VGND VPWR VPWR _124_\[12\] sky130_fd_sc_hd__dfxtp_1
X_13799_ clknet_leaf_61_clk _01018_ VGND VGND VPWR VPWR _128_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12819_ _06453_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__clkbuf_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08010_ _02540_ _02543_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__xor2_1
XFILLER_30_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09961_ _142_\[18\] _04340_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08912_ _03310_ _03311_ _03331_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__and3_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09892_ _142_\[15\] _04274_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__and2_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _228_\[13\] _231_\[13\] _03264_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__o21a_1
X_08774_ _02017_ _03197_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__xor2_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07725_ _02244_ _02246_ _02267_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07656_ _01412_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__clkbuf_4
XFILLER_53_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06607_ _01208_ _01306_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__or2_1
X_07587_ _182_\[15\] _01654_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__nor2_1
XFILLER_43_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06538_ _01207_ _392_\[4\] _01208_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__or3b_4
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09326_ _03698_ _03703_ _03699_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__a21bo_1
X_09257_ _03665_ _03666_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__xnor2_2
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08208_ _164_\[5\] _02701_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__or2_1
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09188_ _170_\[24\] _02849_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__nand2_1
XFILLER_134_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08139_ _167_\[17\] _02652_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__or2_1
XFILLER_107_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11150_ _05227_ _05240_ _05241_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__a21o_1
X_10101_ _04085_ _04177_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__nand2_1
XFILLER_134_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11081_ _03866_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__inv_2
XFILLER_76_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10032_ _04129_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__buf_2
XFILLER_88_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13722_ clknet_leaf_57_clk _00941_ VGND VGND VPWR VPWR _134_\[26\] sky130_fd_sc_hd__dfxtp_1
X_11983_ _05978_ _05979_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10934_ net38 _05068_ _05096_ _05086_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__a211o_1
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13653_ clknet_leaf_47_clk _00872_ VGND VGND VPWR VPWR _138_\[21\] sky130_fd_sc_hd__dfxtp_1
X_10865_ _164_\[23\] _04983_ _05047_ _04998_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__o211a_1
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ clknet_leaf_45_clk _00803_ VGND VGND VPWR VPWR _142_\[16\] sky130_fd_sc_hd__dfxtp_1
X_12604_ _128_\[27\] _126_\[27\] _06335_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__mux2_1
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12535_ _130_\[26\] _128_\[26\] _06302_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__mux2_1
XFILLER_83_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10796_ _164_\[3\] _04983_ _04997_ _04998_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__o211a_1
XFILLER_145_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12466_ _06268_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11417_ _05470_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__clkbuf_1
X_12397_ _132_\[24\] _134_\[24\] _06230_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__mux2_1
X_11348_ _05408_ _05409_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__nor2_1
XFILLER_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11279_ _05348_ _05349_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__or2b_1
XFILLER_67_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13018_ clknet_leaf_12_clk _00237_ VGND VGND VPWR VPWR _240_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07510_ _01642_ _01827_ _01693_ _02060_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__a211o_1
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08490_ _228_\[2\] _231_\[2\] _02776_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__a21o_1
X_07441_ _01991_ _01993_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__or2_1
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07372_ _01927_ _01899_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__or2_1
XFILLER_50_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09111_ _02323_ _03524_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09042_ _03441_ _03442_ _03456_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__o21ai_1
XFILLER_117_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09944_ _246_\[17\] _01315_ _04129_ _243_\[17\] _01482_ VGND VGND VPWR VPWR _04325_
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09875_ _03910_ _01236_ _04179_ _04258_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__or4_1
XFILLER_98_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08826_ _01354_ _03248_ _01412_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__o21ai_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08757_ _03128_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__inv_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _243_\[19\] _240_\[19\] _01667_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__mux2_4
XFILLER_54_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08688_ _03111_ _03114_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _185_\[17\] _234_\[17\] VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__or2_1
XFILLER_41_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10650_ _173_\[24\] _176_\[24\] _01215_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__mux2_1
XFILLER_139_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09309_ _02486_ _03716_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__xor2_1
XFILLER_139_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10581_ _176_\[1\] net68 _01741_ _04682_ _02711_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__a221o_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12320_ _136_\[20\] _134_\[20\] _06189_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__mux2_1
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12251_ _06155_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11202_ _05264_ _05268_ _05275_ _05272_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__o211a_1
XFILLER_79_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12182_ _06119_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11133_ net11 _05202_ _05193_ _158_\[10\] VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__a22o_1
XFILLER_103_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11064_ _164_\[26\] _01218_ _04648_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__o21a_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10015_ _04356_ _04376_ _04392_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__o21ba_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11966_ _05964_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13705_ clknet_leaf_55_clk _00924_ VGND VGND VPWR VPWR _134_\[9\] sky130_fd_sc_hd__dfxtp_1
X_10917_ _167_\[7\] _05036_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__or2_1
X_13636_ clknet_leaf_53_clk _00855_ VGND VGND VPWR VPWR _138_\[4\] sky130_fd_sc_hd__dfxtp_1
X_11897_ _05901_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10848_ _164_\[18\] _05025_ _05034_ _05035_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__a211o_1
X_13567_ clknet_leaf_68_clk _00786_ VGND VGND VPWR VPWR _149_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10779_ _04682_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__clkbuf_4
X_13498_ clknet_leaf_50_clk _00717_ VGND VGND VPWR VPWR _158_\[16\] sky130_fd_sc_hd__dfxtp_1
X_12518_ _130_\[18\] _128_\[18\] _06291_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__mux2_1
XFILLER_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12449_ _132_\[17\] _130_\[17\] _06258_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__mux2_1
XFILLER_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07990_ _02518_ _02523_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__nor2_1
XFILLER_113_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06941_ _01448_ _01555_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__or2_1
X_09660_ _03884_ _04051_ _03925_ _03930_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__a31o_1
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06872_ _01448_ _01505_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__or2_1
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08611_ _03037_ _03039_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__xnor2_4
X_09591_ _03981_ _03982_ _03985_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__a21bo_1
XFILLER_95_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08542_ _170_\[4\] _02781_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__nand2_1
XFILLER_51_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08473_ _02884_ _02906_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__xnor2_1
X_07424_ _01675_ _01976_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__xnor2_2
XFILLER_23_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07355_ _01877_ _01881_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__or2_1
XFILLER_50_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07286_ _01807_ _01836_ _01843_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__and3_1
XFILLER_136_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09025_ _03419_ _03421_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__nor2_1
XFILLER_117_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09927_ _04275_ _04297_ _04307_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__or3b_1
XFILLER_77_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09858_ _04207_ _04219_ _04242_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__o21ba_1
XFILLER_100_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _04155_ _04168_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__nor2_1
XFILLER_100_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08809_ _228_\[12\] _231_\[12\] _03231_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__o21a_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ net31 _05776_ _01368_ _05831_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__a211o_1
XFILLER_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _140_\[20\] _05767_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__xnor2_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_16
X_10702_ _167_\[8\] _04836_ _04931_ _04914_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__a211o_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _05705_ _05706_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__nand2_1
XFILLER_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10633_ _02237_ _04685_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__or2_1
XFILLER_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13421_ clknet_leaf_1_clk _00640_ VGND VGND VPWR VPWR _164_\[7\] sky130_fd_sc_hd__dfxtp_2
X_10564_ _176_\[28\] _04833_ _04806_ _04837_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__o211a_1
XFILLER_6_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13352_ clknet_leaf_0_clk _00571_ VGND VGND VPWR VPWR _170_\[2\] sky130_fd_sc_hd__dfxtp_1
X_12303_ _136_\[12\] _134_\[12\] _06178_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__mux2_1
X_10495_ _04766_ _04788_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__or2_1
X_13283_ clknet_leaf_3_clk _00502_ VGND VGND VPWR VPWR _179_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12234_ _138_\[11\] _136_\[11\] _06145_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__mux2_1
XFILLER_135_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12165_ _06110_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__clkbuf_1
X_11116_ net7 _05215_ _05195_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__mux2_1
XFILLER_68_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12096_ _06074_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11047_ _164_\[19\] _04872_ _04633_ _05169_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__o211a_1
XFILLER_91_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 din[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12998_ clknet_leaf_22_clk _00217_ VGND VGND VPWR VPWR _240_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11949_ _152_\[19\] _05933_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_71_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_51_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13619_ clknet_leaf_46_clk _00838_ VGND VGND VPWR VPWR _140_\[19\] sky130_fd_sc_hd__dfxtp_2
X_07140_ _01670_ _01705_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__or2_1
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07071_ _240_\[14\] _01649_ _01607_ _01652_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__a211o_1
XFILLER_99_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09712_ _03886_ _04025_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__or2_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07973_ _185_\[28\] _234_\[28\] VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__or2_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06924_ _240_\[8\] _01526_ _01510_ _01543_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__o211a_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09643_ _04030_ _04034_ _04024_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__o21ai_1
X_06855_ _243_\[21\] _01474_ _01461_ _01493_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__o211a_1
X_09574_ _03943_ _03968_ _03969_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__or3_1
XFILLER_83_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06786_ _179_\[4\] _01299_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__or2_1
X_08525_ _01789_ _02956_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__xnor2_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_62_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_51_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08456_ _01727_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__inv_2
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07407_ _01959_ _01960_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08387_ _02833_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07338_ _01645_ _237_\[0\] VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07269_ _182_\[5\] _01620_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__or2_1
XFILLER_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10280_ _04630_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09008_ _03422_ _03424_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13970_ clknet_leaf_96_clk _01189_ VGND VGND VPWR VPWR _118_\[18\] sky130_fd_sc_hd__dfxtp_2
X_12921_ clknet_leaf_73_clk _00145_ VGND VGND VPWR VPWR _116_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12852_ _06470_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_53_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_16
X_11803_ _05815_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__inv_2
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12783_ _122_\[16\] _120_\[16\] _06434_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__mux2_1
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _05745_ _05752_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__xor2_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11665_ _149_\[25\] _05279_ _05690_ _05691_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__o22a_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10616_ _176_\[12\] _04872_ _04633_ _04873_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__o211a_1
Xclkbuf_4_6_0_clk clknet_3_3_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_13404_ clknet_leaf_126_clk _00623_ VGND VGND VPWR VPWR _167_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11596_ _116_\[18\] _05628_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__or2_1
XFILLER_128_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13335_ clknet_leaf_8_clk _00554_ VGND VGND VPWR VPWR _173_\[17\] sky130_fd_sc_hd__dfxtp_1
X_10547_ _173_\[23\] _04818_ _04825_ _04823_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__o211a_1
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13266_ clknet_leaf_26_clk _00485_ VGND VGND VPWR VPWR _179_\[12\] sky130_fd_sc_hd__dfxtp_1
X_10478_ _01418_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__buf_2
X_12217_ _138_\[3\] _136_\[3\] _06134_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__mux2_1
X_13197_ clknet_leaf_34_clk _00416_ VGND VGND VPWR VPWR _185_\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_111_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12148_ _140_\[2\] _138_\[2\] _06101_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__mux2_1
XFILLER_96_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12079_ _06065_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06640_ _01246_ _01250_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__nor2_1
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06571_ _01279_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09290_ _170_\[26\] _02855_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__nand2_1
X_08310_ _01406_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__buf_2
XANTENNA_14 _164_\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08241_ _231_\[14\] _02690_ _02712_ _02725_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__a211o_1
XANTENNA_47 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_58 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 _02237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08172_ _02625_ _02675_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__or2_1
X_07123_ _240_\[26\] _01660_ _01653_ _01692_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__o211a_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07054_ _01427_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__buf_2
XFILLER_133_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07956_ _02453_ _02454_ _02491_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__a21oi_1
X_06907_ _176_\[3\] _01531_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__or2_1
XFILLER_56_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07887_ _02422_ _02423_ _02424_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__nand3_1
XFILLER_28_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09626_ _03996_ _04018_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__nand2_1
X_06838_ _01480_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__buf_2
XFILLER_56_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09557_ _01240_ _03927_ _03952_ _01283_ _195_\[4\] VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__a221o_1
XFILLER_55_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06769_ _01427_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__buf_4
X_09488_ _03885_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_35_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
X_08508_ _170_\[3\] _225_\[3\] VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__or2_1
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08439_ _02811_ _02776_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11450_ _05497_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11381_ _01361_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__clkbuf_4
X_10401_ _01225_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__buf_2
XFILLER_109_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10332_ _179_\[25\] _04658_ _04672_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__a21o_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13120_ clknet_leaf_117_clk _00339_ VGND VGND VPWR VPWR _228_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13051_ clknet_leaf_85_clk _00270_ VGND VGND VPWR VPWR _237_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12002_ _152_\[25\] _05995_ _05996_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__and3_1
X_10263_ _04628_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__buf_4
XFILLER_132_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10194_ _04561_ _04563_ _01233_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__mux2_1
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13953_ clknet_leaf_70_clk _01172_ VGND VGND VPWR VPWR _118_\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_19_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13884_ clknet_leaf_72_clk _01103_ VGND VGND VPWR VPWR _124_\[28\] sky130_fd_sc_hd__dfxtp_1
X_12904_ clknet_leaf_93_clk _00128_ VGND VGND VPWR VPWR _116_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _06461_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _122_\[8\] _120_\[8\] _06423_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__mux2_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _06389_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__clkbuf_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _118_\[17\] _116_\[31\] VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__xor2_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 din[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
X_11648_ _118_\[27\] _118_\[31\] VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11579_ _05612_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__xor2_1
Xinput34 rst VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_4
Xinput23 din[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
XFILLER_115_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13318_ clknet_leaf_23_clk _00537_ VGND VGND VPWR VPWR _173_\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_10_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13249_ clknet_leaf_7_clk _00468_ VGND VGND VPWR VPWR _182_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07810_ _02289_ _02296_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__nand2_1
X_08790_ _03179_ _03213_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__nor2_1
XFILLER_84_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07741_ _182_\[17\] _01661_ _02227_ _02228_ _02235_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__o2111ai_1
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07672_ _02215_ _02216_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06623_ _01247_ _01272_ _01307_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__nand3_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09411_ _02835_ _03815_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06554_ _158_\[17\] _158_\[16\] _01262_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_17_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_80_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09342_ _02506_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__xor2_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09273_ _02460_ _03681_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08224_ _228_\[9\] _02698_ _02679_ _02713_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__o211a_1
XFILLER_107_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08155_ _01435_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07106_ _01670_ _01679_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__or2_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08086_ _01670_ _02614_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__or2_1
XFILLER_134_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07037_ _237_\[7\] VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__buf_6
XFILLER_88_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08988_ _03372_ _03375_ _03371_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__o21ai_2
X_07939_ _02473_ _02475_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__xnor2_2
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10950_ _01225_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09609_ _03890_ _03896_ _03927_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__a31oi_1
XFILLER_113_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10881_ _164_\[28\] _05025_ _05058_ _05035_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__a211o_1
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12620_ _06349_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12551_ _06200_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__buf_4
XFILLER_138_830 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12482_ _130_\[1\] _128_\[1\] _06269_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__mux2_1
X_11502_ _149_\[8\] _05545_ _05533_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__mux2_1
XFILLER_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11433_ _05483_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11364_ _05421_ _05423_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11295_ _05342_ _05344_ _05349_ _05363_ _05348_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__a311o_1
X_10315_ _04633_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13103_ clknet_leaf_117_clk _00322_ VGND VGND VPWR VPWR _231_\[15\] sky130_fd_sc_hd__dfxtp_1
X_10246_ _142_\[30\] _04601_ _04602_ _04600_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__a22o_1
XFILLER_106_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13034_ clknet_leaf_45_clk _00253_ VGND VGND VPWR VPWR _237_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10177_ _04515_ _04524_ _04547_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__nor3b_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13936_ clknet_leaf_96_clk _01155_ VGND VGND VPWR VPWR _120_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13867_ clknet_leaf_95_clk _01086_ VGND VGND VPWR VPWR _124_\[11\] sky130_fd_sc_hd__dfxtp_1
X_13798_ clknet_leaf_60_clk _01017_ VGND VGND VPWR VPWR _128_\[6\] sky130_fd_sc_hd__dfxtp_1
X_12818_ _118_\[1\] _120_\[1\] _06451_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__mux2_1
XFILLER_43_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12749_ _122_\[0\] _120_\[0\] _06412_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__mux2_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09960_ _246_\[18\] _01315_ _04129_ _243_\[18\] _01486_ VGND VGND VPWR VPWR _04340_
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_6_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08911_ _03329_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__nor2_1
XFILLER_112_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09891_ _246_\[15\] _01314_ _04129_ _243_\[15\] _01475_ VGND VGND VPWR VPWR _04274_
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _228_\[13\] _231_\[13\] _02811_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__a21o_1
XFILLER_85_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08773_ _03194_ _03196_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__xnor2_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07724_ _02265_ _02266_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__nand2_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07655_ _02197_ _02199_ _02200_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__a21o_1
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06606_ _01308_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__inv_2
XFILLER_25_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07586_ _02131_ _02133_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__xnor2_1
X_06537_ _01245_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__buf_2
X_09325_ _170_\[27\] _02858_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__xnor2_2
XFILLER_139_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09256_ _03600_ _03606_ _03599_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__o21a_1
X_08207_ _01339_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__clkbuf_2
XFILLER_107_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09187_ _170_\[24\] _02849_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__or2_1
XFILLER_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08138_ _01339_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__clkbuf_2
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08069_ _02598_ _02600_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__xnor2_1
X_10100_ _04472_ _04473_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__or2_1
XFILLER_108_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11080_ _03866_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__inv_2
X_10031_ _185_\[20\] _03870_ _04175_ _04408_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__o211a_1
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13721_ clknet_leaf_56_clk _00940_ VGND VGND VPWR VPWR _134_\[25\] sky130_fd_sc_hd__dfxtp_1
X_11982_ _05967_ _05970_ _05966_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__a21bo_1
XFILLER_91_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10933_ _164_\[11\] _05059_ _05094_ _05095_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__o211a_1
XFILLER_32_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13652_ clknet_leaf_48_clk _00871_ VGND VGND VPWR VPWR _138_\[20\] sky130_fd_sc_hd__dfxtp_1
X_10864_ _05028_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__or2_1
XFILLER_140_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13583_ clknet_leaf_45_clk _00802_ VGND VGND VPWR VPWR _142_\[15\] sky130_fd_sc_hd__dfxtp_1
X_12603_ _06340_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__clkbuf_1
X_10795_ _01424_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__clkbuf_4
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12534_ _06304_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12465_ _132_\[25\] _130_\[25\] _06258_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__mux2_1
X_11416_ _152_\[30\] _05469_ _05439_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__mux2_1
X_12396_ _06232_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11347_ _149_\[22\] _132_\[22\] VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__and2_1
XFILLER_98_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11278_ _149_\[13\] _132_\[13\] VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__nand2_1
X_10229_ _03950_ _04363_ _03890_ _04437_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__o211a_1
X_13017_ clknet_leaf_14_clk _00236_ VGND VGND VPWR VPWR _240_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13919_ clknet_leaf_69_clk _01138_ VGND VGND VPWR VPWR _122_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07440_ _01944_ _01992_ _01962_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07371_ _01896_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__inv_2
X_09110_ _03522_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__nand2_1
X_09041_ _03441_ _03442_ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__nor3_1
XFILLER_30_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09943_ _04315_ _04317_ _04323_ _04210_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__o22a_1
X_09874_ _04002_ _03888_ _03929_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__and3_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _03245_ _03247_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08756_ _03179_ _03180_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__or2_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07707_ _02248_ _02250_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__xnor2_1
X_08687_ _03112_ _03113_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__nor2_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _01698_ _02183_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__xnor2_2
XFILLER_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07569_ _02116_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__inv_2
XFILLER_110_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09308_ _03714_ _03715_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__nand2_1
XFILLER_139_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10580_ _04848_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__clkbuf_4
XFILLER_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09239_ _03647_ _03648_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__and2_1
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12250_ _138_\[19\] _136_\[19\] _06145_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__mux2_1
X_11201_ _05280_ _05281_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__or2b_1
XFILLER_123_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12181_ _140_\[18\] _138_\[18\] _06112_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__mux2_1
X_11132_ _158_\[10\] _01258_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11063_ _03667_ _05110_ _05179_ _01436_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__a211o_1
X_10014_ _04390_ _04391_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__or2b_1
XFILLER_89_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11965_ _142_\[21\] _05963_ _05893_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__mux2_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13704_ clknet_leaf_54_clk _00923_ VGND VGND VPWR VPWR _134_\[8\] sky130_fd_sc_hd__dfxtp_1
X_10916_ net64 _05048_ _05083_ _05067_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__o211a_1
X_13635_ clknet_leaf_53_clk _00854_ VGND VGND VPWR VPWR _138_\[3\] sky130_fd_sc_hd__dfxtp_1
X_11896_ _142_\[15\] _05900_ _05893_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__mux2_1
XFILLER_72_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10847_ _01418_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__clkbuf_4
XFILLER_20_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13566_ clknet_leaf_75_clk _00785_ VGND VGND VPWR VPWR _149_\[30\] sky130_fd_sc_hd__dfxtp_1
X_10778_ _167_\[30\] _04983_ _04985_ _04939_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__o211a_1
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13497_ clknet_leaf_41_clk _00716_ VGND VGND VPWR VPWR _158_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12517_ _06295_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12448_ _06259_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12379_ _06223_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06940_ _176_\[13\] _240_\[13\] _01449_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__mux2_1
XFILLER_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06871_ _179_\[26\] _243_\[26\] _01449_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__mux2_1
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08610_ _03004_ _03007_ _03038_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__o21ai_2
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09590_ _03876_ _03928_ _03984_ _03880_ _195_\[4\] VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__a221o_1
XFILLER_82_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08541_ _170_\[4\] _02781_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__nor2_1
XFILLER_35_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08472_ _170_\[1\] _02772_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__xor2_2
XFILLER_35_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07423_ _01657_ _01612_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07354_ _01910_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__inv_2
XFILLER_108_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07285_ _01807_ _01836_ _01843_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__a21oi_1
XFILLER_136_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09024_ _02827_ _01426_ _03379_ _03440_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__o211a_1
XFILLER_117_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09926_ _04275_ _04297_ _04307_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__o21bai_2
XFILLER_86_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09857_ _04240_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__or2_1
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _02833_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__buf_2
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08808_ _228_\[12\] _231_\[12\] _02807_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__a21o_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _01985_ _03163_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _140_\[22\] _140_\[13\] VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _170_\[8\] _04833_ _04922_ _04930_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__o211a_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11681_ _116_\[27\] _05704_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__or2_1
XFILLER_139_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10632_ _04855_ _04882_ _04883_ _04839_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__a211o_1
X_13420_ clknet_leaf_113_clk _00639_ VGND VGND VPWR VPWR _164_\[6\] sky130_fd_sc_hd__dfxtp_1
X_10563_ _179_\[28\] _04799_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__or2_1
X_13351_ clknet_leaf_2_clk _00570_ VGND VGND VPWR VPWR _170_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12302_ _06182_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10494_ _176_\[8\] _179_\[8\] _04743_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__mux2_1
X_13282_ clknet_leaf_8_clk _00501_ VGND VGND VPWR VPWR _179_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12233_ _06146_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12164_ _140_\[10\] _138_\[10\] _06101_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__mux2_1
X_12095_ _140_\[9\] _142_\[9\] _06068_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__mux2_1
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11115_ _01256_ _05214_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__nand2_1
XFILLER_122_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11046_ _03464_ _04681_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__nand2_1
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12997_ clknet_leaf_19_clk _00216_ VGND VGND VPWR VPWR _240_\[5\] sky130_fd_sc_hd__dfxtp_1
X_11948_ _05925_ _05947_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__or2_1
XFILLER_60_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11879_ _140_\[24\] _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__xnor2_2
X_13618_ clknet_leaf_49_clk _00837_ VGND VGND VPWR VPWR _140_\[18\] sky130_fd_sc_hd__dfxtp_2
X_13549_ clknet_leaf_87_clk _00768_ VGND VGND VPWR VPWR _149_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07070_ _01650_ _01639_ _01609_ _01651_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__o211a_1
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09711_ _142_\[7\] _04073_ _04100_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07972_ _185_\[28\] _234_\[28\] VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__nand2_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06923_ _176_\[8\] _01531_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__or2_1
XFILLER_68_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09642_ _04024_ _04030_ _04034_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__or3_1
X_06854_ _179_\[21\] _01301_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__or2_1
XFILLER_95_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09573_ _03948_ _03949_ _03967_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__nor3_1
X_06785_ _246_\[3\] _01407_ _01436_ _01441_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__a211o_1
XFILLER_83_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08524_ _02953_ _02955_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__xor2_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08455_ _02880_ _02882_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__and2b_1
XFILLER_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07406_ _243_\[9\] _240_\[9\] _01632_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__mux2_2
XFILLER_51_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08386_ _01423_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__buf_6
X_07337_ _01867_ _01868_ _01869_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__nand3_1
XFILLER_109_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07268_ _01406_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07199_ _01759_ _01760_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__xnor2_1
X_09007_ _228_\[18\] _231_\[18\] _03423_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__o21a_1
XFILLER_104_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09909_ _04289_ _04291_ _03945_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12920_ clknet_leaf_73_clk _00144_ VGND VGND VPWR VPWR _116_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12851_ _118_\[17\] _120_\[17\] _06462_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__mux2_1
X_11802_ _152_\[7\] _05813_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__nor2_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _01392_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__buf_4
XFILLER_14_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _152_\[1\] _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__xnor2_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11664_ _05688_ _05689_ _05263_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__o21ai_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10615_ _02058_ _04872_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__nand2_1
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13403_ clknet_leaf_125_clk _00622_ VGND VGND VPWR VPWR _167_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11595_ _116_\[18\] _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__nand2_1
X_13334_ clknet_leaf_5_clk _00553_ VGND VGND VPWR VPWR _173_\[16\] sky130_fd_sc_hd__dfxtp_2
X_10546_ _04809_ _04824_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__or2_1
XFILLER_10_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13265_ clknet_leaf_25_clk _00484_ VGND VGND VPWR VPWR _179_\[11\] sky130_fd_sc_hd__dfxtp_1
X_10477_ _176_\[3\] _04771_ _04751_ _04775_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__o211a_1
XFILLER_51_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12216_ _06137_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__clkbuf_1
X_13196_ clknet_leaf_34_clk _00415_ VGND VGND VPWR VPWR _185_\[6\] sky130_fd_sc_hd__dfxtp_2
X_12147_ _01393_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__clkbuf_4
XFILLER_123_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12078_ _140_\[1\] _142_\[1\] _06005_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__mux2_1
XFILLER_111_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11029_ _164_\[13\] _01217_ _04627_ net40 _05157_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__o221a_1
XFILLER_37_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06570_ _195_\[1\] VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__buf_2
XFILLER_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08240_ _228_\[14\] _02698_ _02723_ _02724_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__o211a_1
XFILLER_33_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_26 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08171_ _167_\[27\] _231_\[27\] _02626_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__mux2_1
XANTENNA_15 _164_\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_59 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07122_ _01670_ _01691_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__or2_1
XFILLER_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07053_ _237_\[11\] VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__buf_4
XFILLER_114_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07955_ _02489_ _02490_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__nand2_1
XFILLER_101_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06906_ _01339_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__clkbuf_2
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09625_ _03996_ _04018_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__or2_1
XFILLER_83_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07886_ _185_\[25\] _234_\[25\] VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__nand2_1
XFILLER_28_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06837_ _01423_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__buf_4
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09556_ _03951_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__buf_2
XFILLER_71_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06768_ _01408_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__buf_4
X_09487_ _01277_ _01282_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__and2_1
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06699_ _118_\[14\] _116_\[14\] _01381_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__mux2_1
X_08507_ _02939_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__clkbuf_1
X_08438_ _228_\[31\] _02838_ _02861_ _02873_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__a211o_1
XFILLER_11_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08369_ _225_\[16\] VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__clkbuf_4
X_11380_ _05435_ _05437_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__xnor2_1
X_10400_ _176_\[13\] _04691_ _04720_ _04677_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__o211a_1
X_10331_ _182_\[25\] _04654_ _04671_ _04650_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__a31o_1
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13050_ clknet_leaf_108_clk _00269_ VGND VGND VPWR VPWR _237_\[26\] sky130_fd_sc_hd__dfxtp_1
X_10262_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__clkbuf_4
X_12001_ _140_\[10\] _140_\[12\] VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__nand2_1
XFILLER_3_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10193_ _01239_ _03890_ _03888_ _03938_ _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__a41o_1
XFILLER_127_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13952_ clknet_leaf_70_clk _01171_ VGND VGND VPWR VPWR _118_\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12903_ clknet_leaf_91_clk _00127_ VGND VGND VPWR VPWR _116_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13883_ clknet_leaf_89_clk _01102_ VGND VGND VPWR VPWR _124_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _118_\[9\] _120_\[9\] _06451_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__mux2_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _06425_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__clkbuf_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _05725_ _05731_ _05733_ _05732_ _116_\[30\] VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__a32o_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12696_ _124_\[7\] _122_\[7\] _06379_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__mux2_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11647_ _05675_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__clkbuf_1
Xinput13 din[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
Xinput24 din[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput35 src_ready VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_6
X_11578_ _05595_ _05597_ _05604_ _05613_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__o31a_1
XFILLER_7_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10529_ _176_\[18\] _04771_ _04806_ _04812_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__o211a_1
X_13317_ clknet_leaf_10_clk _00536_ VGND VGND VPWR VPWR _176_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13248_ clknet_leaf_5_clk _00467_ VGND VGND VPWR VPWR _182_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13179_ clknet_leaf_102_clk _00398_ VGND VGND VPWR VPWR _225_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07740_ _182_\[18\] _01664_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__nand2_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07671_ _243_\[18\] _240_\[18\] _01664_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__mux2_4
XFILLER_53_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06622_ _01207_ _01310_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__or2_2
XFILLER_53_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09410_ _02804_ _02768_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__xnor2_1
X_06553_ _158_\[15\] _01261_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__or2_1
X_09341_ _03746_ _03747_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__nand2_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09272_ _03679_ _03680_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__and2_1
XFILLER_21_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08223_ _164_\[9\] _02701_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__or2_1
XFILLER_119_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08154_ _234_\[21\] _02659_ _02636_ _02663_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__o211a_1
XFILLER_107_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07105_ _173_\[22\] _01678_ _01672_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__mux2_1
X_08085_ _167_\[2\] _231_\[2\] _01672_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__mux2_1
X_07036_ _240_\[6\] _01601_ _01598_ _01625_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__o211a_1
XFILLER_106_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_clk clknet_3_2_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08987_ _03403_ _03404_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__nand2_1
XFILLER_102_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07938_ _02441_ _02444_ _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__a21o_1
XFILLER_29_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07869_ _182_\[20\] _01671_ _02285_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__o21ba_1
X_09608_ _03879_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__buf_2
XFILLER_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10880_ _167_\[28\] _05022_ _05043_ _05057_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__o211a_1
X_09539_ _01277_ _03877_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__and2_1
XFILLER_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12550_ _06312_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12481_ _06276_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__clkbuf_1
X_11501_ _05539_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__xor2_1
XFILLER_8_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11432_ _149_\[1\] _05482_ _05439_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__mux2_1
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11363_ _05409_ _05414_ _05422_ _05416_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__o31a_1
XFILLER_98_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13102_ clknet_leaf_116_clk _00321_ VGND VGND VPWR VPWR _231_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11294_ _05356_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__inv_2
X_10314_ _182_\[17\] _04634_ _04662_ _04649_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__o211a_1
X_13033_ clknet_leaf_42_clk _00252_ VGND VGND VPWR VPWR _237_\[9\] sky130_fd_sc_hd__dfxtp_1
X_10245_ _01353_ _04611_ _01521_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__a21oi_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10176_ _04539_ _04546_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13935_ clknet_leaf_97_clk _01154_ VGND VGND VPWR VPWR _120_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13866_ clknet_leaf_97_clk _01085_ VGND VGND VPWR VPWR _124_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12817_ _06452_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__clkbuf_1
X_13797_ clknet_leaf_63_clk _01016_ VGND VGND VPWR VPWR _128_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12748_ _06416_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__clkbuf_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ _06380_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09890_ _185_\[14\] _04150_ _04175_ _04273_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__o211a_1
X_08910_ _03288_ _03312_ _03328_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__o21a_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08841_ _03260_ _03262_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__xnor2_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08772_ _02006_ _03159_ _03195_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__o21a_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07723_ _02263_ _02264_ _02262_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__a21o_1
XFILLER_93_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07654_ _02197_ _02199_ _01519_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06605_ _01297_ _01307_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__nor2_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07585_ _02101_ _02104_ _02132_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__a21bo_1
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06536_ _392_\[3\] _392_\[2\] VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__or2b_1
X_09324_ _03689_ _03696_ _03730_ _01408_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__a31o_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09255_ _03663_ _03664_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__and2_1
X_08206_ _231_\[4\] _02690_ _02664_ _02700_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__a211o_1
X_09186_ _02846_ _01426_ _03379_ _03597_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__o211a_1
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08137_ _234_\[16\] _02646_ _02629_ _02651_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__a211o_1
X_08068_ _234_\[31\] _02599_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07019_ _237_\[3\] VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__buf_4
XFILLER_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10030_ _04406_ _04407_ _03945_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__a21o_1
XFILLER_88_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11981_ _05976_ _05977_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__or2b_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13720_ clknet_leaf_67_clk _00939_ VGND VGND VPWR VPWR _134_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10932_ _167_\[11\] _05089_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__or2_1
XFILLER_140_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13651_ clknet_leaf_77_clk _00870_ VGND VGND VPWR VPWR _138_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10863_ _167_\[23\] _170_\[23\] _04995_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__mux2_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13582_ clknet_leaf_45_clk _00801_ VGND VGND VPWR VPWR _142_\[14\] sky130_fd_sc_hd__dfxtp_1
X_12602_ _128_\[26\] _126_\[26\] _06335_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__mux2_1
X_10794_ _04971_ _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__or2_1
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12533_ _130_\[25\] _128_\[25\] _06302_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__mux2_1
XFILLER_8_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12464_ _06267_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11415_ _05466_ _05468_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__xnor2_1
X_12395_ _132_\[23\] _134_\[23\] _06230_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__mux2_1
X_11346_ _149_\[22\] _132_\[22\] VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__nor2_1
XFILLER_4_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11277_ _149_\[13\] _132_\[13\] VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__nor2_1
X_13016_ clknet_leaf_14_clk _00235_ VGND VGND VPWR VPWR _240_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10228_ _04164_ _04386_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__nor2_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10159_ _04451_ _04452_ _04489_ _04490_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__o311ai_4
XFILLER_79_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13918_ clknet_leaf_68_clk _01137_ VGND VGND VPWR VPWR _122_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13849_ clknet_leaf_90_clk _01068_ VGND VGND VPWR VPWR _126_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07370_ _01903_ _01906_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__and2b_1
XFILLER_31_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09040_ _03453_ _03455_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09942_ _04319_ _04322_ _01237_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__mux2_1
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09873_ _03871_ _04078_ _04132_ _04058_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__or4_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _03210_ _03246_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__nor2_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08755_ _170_\[10\] _02801_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__nor2_1
X_07706_ _02249_ _02211_ _02210_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__o21a_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08686_ _228_\[8\] _231_\[8\] _02794_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__a21oi_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07637_ _01681_ _01635_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07568_ _01690_ _02115_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__xnor2_1
X_06519_ _01227_ _01219_ _01228_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__and3_1
X_09307_ _185_\[27\] _03713_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__or2_1
X_07499_ _02014_ _02036_ _02049_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__o21a_1
X_09238_ _03640_ _03642_ _03646_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__nand3_1
X_09169_ _02371_ _03580_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11200_ _149_\[3\] _132_\[3\] VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__nand2_1
XFILLER_119_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12180_ _06118_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11131_ _05191_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11062_ net53 _01226_ _04865_ _05178_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__o211a_1
XFILLER_1_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10013_ _04381_ _04389_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__nand2_1
XFILLER_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11964_ net14 _05962_ _05852_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__mux2_1
X_13703_ clknet_leaf_59_clk _00922_ VGND VGND VPWR VPWR _134_\[7\] sky130_fd_sc_hd__dfxtp_1
X_11895_ net7 _05899_ _05852_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__mux2_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10915_ _05079_ _05082_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__or2_1
XFILLER_17_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13634_ clknet_leaf_54_clk _00853_ VGND VGND VPWR VPWR _138_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10846_ _167_\[18\] _05022_ _05009_ _05033_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__o211a_1
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13565_ clknet_leaf_76_clk _00784_ VGND VGND VPWR VPWR _149_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10777_ _04971_ _04984_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__or2_1
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13496_ clknet_leaf_41_clk _00715_ VGND VGND VPWR VPWR _158_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12516_ _130_\[17\] _128_\[17\] _06291_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__mux2_1
XFILLER_145_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12447_ _132_\[16\] _130_\[16\] _06258_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__mux2_1
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12378_ _132_\[15\] _134_\[15\] _06219_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__mux2_1
XFILLER_114_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11329_ _05393_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06870_ _246_\[25\] _01496_ _01460_ _01504_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__a211o_1
XFILLER_94_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08540_ _225_\[3\] _02845_ _02834_ _02971_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__o211a_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08471_ _02889_ _02903_ _01518_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__o21ai_1
X_07422_ _01974_ _01955_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__or2_1
XFILLER_51_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07353_ _01908_ _01909_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__or2b_1
X_07284_ _01841_ _01842_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__nand2_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09023_ _03432_ _03433_ _03439_ _02355_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__a211o_1
XFILLER_144_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09925_ _04299_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09856_ _04229_ _04239_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__and2_1
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08807_ _03228_ _03229_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__or2b_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _185_\[10\] _04150_ _03919_ _04174_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__o211a_1
XFILLER_100_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06999_ _01568_ _01596_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__or2_1
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _03160_ _03162_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__xor2_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _03070_ _03085_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__nor2_1
XFILLER_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _173_\[8\] _04917_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__or2_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _116_\[27\] _05704_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__nand2_1
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10631_ _02230_ _04631_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__nor2_1
XFILLER_10_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13350_ clknet_leaf_0_clk _00569_ VGND VGND VPWR VPWR _170_\[0\] sky130_fd_sc_hd__dfxtp_2
X_10562_ _04682_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__clkbuf_4
X_12301_ _136_\[11\] _134_\[11\] _06178_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__mux2_1
X_13281_ clknet_leaf_7_clk _00500_ VGND VGND VPWR VPWR _179_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12232_ _138_\[10\] _136_\[10\] _06145_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__mux2_1
X_10493_ _173_\[7\] _04774_ _04787_ _04777_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__a211o_1
XFILLER_6_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12163_ _06109_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12094_ _06073_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11114_ _158_\[6\] _01255_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__nand2_1
XFILLER_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11045_ _03438_ _04861_ _05168_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__a21boi_1
XFILLER_76_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12996_ clknet_leaf_20_clk _00215_ VGND VGND VPWR VPWR _240_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11947_ _05924_ _05936_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__or2_1
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11878_ _140_\[31\] _140_\[1\] VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__xnor2_2
XFILLER_60_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13617_ clknet_leaf_45_clk _00836_ VGND VGND VPWR VPWR _140_\[17\] sky130_fd_sc_hd__dfxtp_2
X_10829_ _164_\[13\] _04986_ _05021_ _05001_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__a211o_1
X_13548_ clknet_leaf_84_clk _00767_ VGND VGND VPWR VPWR _149_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13479_ clknet_leaf_28_clk _00698_ _00112_ VGND VGND VPWR VPWR _190_\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07971_ _01675_ _02505_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__xnor2_4
XFILLER_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09710_ _04074_ _04091_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__nor2_1
XFILLER_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06922_ _243_\[7\] _01536_ _01509_ _01542_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__a211o_1
XFILLER_68_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09641_ _03937_ _03959_ _04033_ _03871_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__a211oi_1
X_06853_ _246_\[20\] _01485_ _01481_ _01492_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__o211a_1
XFILLER_68_787 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09572_ _03948_ _03949_ _03967_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__o21a_1
X_06784_ _243_\[3\] _01438_ _01439_ _01440_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__o211a_1
XFILLER_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08523_ _02911_ _02914_ _02954_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__o21a_1
XFILLER_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08454_ _02768_ _02838_ _02861_ _02888_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__a211o_1
X_07405_ _01957_ _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__or2_1
XFILLER_51_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08385_ _228_\[19\] _02771_ _02765_ _02832_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__o211a_1
XFILLER_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07336_ _01874_ _01875_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__or2b_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07267_ _01616_ _01649_ _01693_ _01826_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__a211o_1
X_09006_ _228_\[18\] _231_\[18\] _02827_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__a21o_1
XFILLER_145_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07198_ _01727_ _01730_ _01728_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09908_ _04266_ _04270_ _04290_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__o21ai_1
XFILLER_76_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09839_ _04205_ _04224_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__or2_1
XFILLER_58_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12850_ _06469_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__clkbuf_1
X_11801_ _152_\[7\] _05813_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__nand2_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12781_ _06433_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _140_\[20\] _05750_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__xnor2_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11663_ _05688_ _05689_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__and2_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10614_ _04636_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__buf_4
X_13402_ clknet_leaf_130_clk _00621_ VGND VGND VPWR VPWR _167_\[20\] sky130_fd_sc_hd__dfxtp_2
X_11594_ _118_\[4\] _05627_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__xnor2_1
X_13333_ clknet_leaf_23_clk _00552_ VGND VGND VPWR VPWR _173_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10545_ _176_\[23\] _179_\[23\] _04790_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__mux2_1
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_130_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_130_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13264_ clknet_leaf_27_clk _00483_ VGND VGND VPWR VPWR _179_\[10\] sky130_fd_sc_hd__dfxtp_1
X_10476_ _179_\[3\] _04746_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__or2_1
XFILLER_6_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12215_ _138_\[2\] _136_\[2\] _06134_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__mux2_1
X_13195_ clknet_leaf_34_clk _00414_ VGND VGND VPWR VPWR _185_\[5\] sky130_fd_sc_hd__dfxtp_4
XFILLER_6_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12146_ _06100_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12077_ _06064_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11028_ _03275_ _04636_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__nand2_1
XFILLER_37_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12979_ clknet_leaf_23_clk _00198_ VGND VGND VPWR VPWR _243_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_27 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08170_ _234_\[26\] _02646_ _02664_ _02674_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__a211o_1
XFILLER_20_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_16 _164_\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_49 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07121_ _173_\[26\] _01690_ _01672_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__mux2_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07052_ _240_\[10\] _01601_ _01598_ _01637_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__o211a_1
XFILLER_99_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07954_ _02487_ _02488_ _02486_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__a21o_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06905_ _243_\[2\] _01485_ _01481_ _01530_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__o211a_1
X_07885_ _185_\[25\] _234_\[25\] VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__or2_1
XFILLER_28_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09624_ _04015_ _04017_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__xor2_2
X_06836_ _246_\[16\] _01422_ _01425_ _01479_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__o211a_1
XFILLER_83_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09555_ _03879_ _03950_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__and2_1
X_06767_ _01412_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__clkbuf_8
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09486_ _01240_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__buf_2
XFILLER_70_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06698_ _01367_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__buf_4
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08506_ _01710_ _02938_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__or2_1
XFILLER_62_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08437_ _02871_ _01801_ _02824_ _02872_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__o211a_1
XFILLER_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08368_ _228_\[15\] _02775_ _02810_ _02819_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__a211o_1
XFILLER_137_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07319_ _01844_ _01865_ _01876_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_112_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_112_clk sky130_fd_sc_hd__clkbuf_16
X_08299_ _02749_ _02766_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__or2_1
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10330_ _04630_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__clkbuf_4
X_10261_ _04626_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__buf_4
XFILLER_117_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12000_ _140_\[10\] _140_\[12\] VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__or2_1
X_10192_ _04303_ _04233_ _04437_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__o21a_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13951_ clknet_leaf_69_clk _01170_ VGND VGND VPWR VPWR _120_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12902_ clknet_leaf_91_clk _00126_ VGND VGND VPWR VPWR _116_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13882_ clknet_leaf_89_clk _01101_ VGND VGND VPWR VPWR _124_\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12833_ _06460_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _122_\[7\] _120_\[7\] _06423_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__mux2_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _05734_ _05736_ _149_\[30\] _05262_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12695_ _06388_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__clkbuf_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11646_ _149_\[23\] _05674_ _05625_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__mux2_1
Xinput25 din[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
Xinput14 din[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
X_11577_ _05593_ _05603_ _05602_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_103_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_103_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10528_ _179_\[18\] _04799_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__or2_1
X_13316_ clknet_leaf_5_clk _00535_ VGND VGND VPWR VPWR _176_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13247_ clknet_leaf_5_clk _00466_ VGND VGND VPWR VPWR _182_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10459_ _04712_ _04762_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__or2_1
XFILLER_123_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13178_ clknet_leaf_101_clk _00397_ VGND VGND VPWR VPWR _225_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12129_ _140_\[25\] _142_\[25\] _06090_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__mux2_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07670_ _02213_ _02214_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__or2_1
XFILLER_38_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06621_ _01207_ _01208_ _01250_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__or3_2
XFILLER_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06552_ _158_\[13\] _158_\[14\] _01260_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__or3_1
X_09340_ _185_\[28\] _03745_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__or2_1
X_09271_ _03672_ _03674_ _03678_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__nand3_1
X_08222_ _02711_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__clkbuf_4
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08153_ _02625_ _02662_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__or2_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08084_ _234_\[1\] _02564_ _02178_ _02613_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__a211o_1
X_07104_ _237_\[22\] VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__buf_6
X_07035_ _01615_ _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__or2_1
XFILLER_115_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08986_ _170_\[17\] _02823_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__or2_1
X_07937_ _182_\[25\] _01687_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__nor2_1
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07868_ _02290_ _02298_ _02350_ _02357_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__or4bb_1
XFILLER_29_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09607_ _03873_ _03893_ _03979_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06819_ _243_\[12\] _01428_ _01466_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07799_ _02308_ _02322_ _02338_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__or3_1
X_09538_ _01277_ _01279_ _01282_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__and3b_2
XFILLER_71_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09469_ _01295_ _01271_ _01272_ _01274_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__o211ai_4
X_11500_ _05542_ _05543_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__nand2_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12480_ _130_\[0\] _128_\[0\] _06269_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__mux2_1
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11431_ _05477_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__xor2_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11362_ _149_\[23\] _132_\[23\] VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__and2_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10313_ _179_\[17\] _04646_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__or2_1
X_13101_ clknet_leaf_116_clk _00320_ VGND VGND VPWR VPWR _231_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11293_ _05360_ _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__or2b_1
XFILLER_133_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13032_ clknet_leaf_42_clk _00251_ VGND VGND VPWR VPWR _237_\[8\] sky130_fd_sc_hd__dfxtp_1
X_10244_ _246_\[31\] _243_\[31\] _01316_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__mux2_1
X_10175_ _04210_ _04541_ _04543_ _04545_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__a31o_1
XFILLER_78_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13934_ clknet_leaf_97_clk _01153_ VGND VGND VPWR VPWR _120_\[14\] sky130_fd_sc_hd__dfxtp_1
X_13865_ clknet_leaf_62_clk _01084_ VGND VGND VPWR VPWR _124_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12816_ _118_\[0\] _120_\[0\] _06451_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__mux2_1
XFILLER_74_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13796_ clknet_leaf_62_clk _01015_ VGND VGND VPWR VPWR _128_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12747_ _124_\[31\] _122_\[31\] _06412_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__mux2_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12678_ _126_\[30\] _124_\[30\] _06379_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__mux2_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11629_ _05646_ _05650_ _05658_ _05352_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__a31o_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08840_ _02048_ _03226_ _03261_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__a21oi_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08771_ _185_\[10\] _03158_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__nand2_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07722_ _02262_ _02263_ _02264_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__nand3_1
XFILLER_93_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07653_ _02198_ _02166_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__and2_1
XFILLER_53_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06604_ _01306_ _01251_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__or2_2
XFILLER_92_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07584_ _02100_ _02098_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__or2b_1
X_09323_ _03689_ _03696_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__a21oi_1
X_06535_ _01243_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__buf_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09254_ _170_\[25\] _02852_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__or2_1
X_08205_ _228_\[4\] _02698_ _02679_ _02699_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__o211a_1
X_09185_ _03591_ _03592_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__a21o_1
XFILLER_119_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08136_ _231_\[16\] _02649_ _02641_ _02650_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__o211a_1
XFILLER_107_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08067_ _02573_ _02576_ _02575_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__a21o_1
XFILLER_115_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07018_ _240_\[2\] _01583_ _01607_ _01611_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__a211o_1
XFILLER_0_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08969_ _02151_ _03345_ _03386_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__o21a_1
X_11980_ _152_\[23\] _05974_ _05975_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__nand3_1
XFILLER_57_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10931_ _04685_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__clkbuf_4
XFILLER_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13650_ clknet_leaf_47_clk _00869_ VGND VGND VPWR VPWR _138_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10862_ _164_\[22\] _05025_ _05045_ _05035_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__a211o_1
X_13581_ clknet_leaf_51_clk _00800_ VGND VGND VPWR VPWR _142_\[13\] sky130_fd_sc_hd__dfxtp_1
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _06339_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10793_ _167_\[3\] _170_\[3\] _04995_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__mux2_1
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ _06303_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12463_ _132_\[24\] _130_\[24\] _06258_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__mux2_1
XFILLER_40_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11414_ _05467_ _05460_ _05458_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__o21ai_1
XFILLER_125_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12394_ _06231_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11345_ _05407_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11276_ _05279_ _05344_ _05346_ _05347_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__a31o_1
XFILLER_4_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10227_ _01239_ _04594_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__nor2_1
X_13015_ clknet_leaf_3_clk _00234_ VGND VGND VPWR VPWR _240_\[23\] sky130_fd_sc_hd__dfxtp_1
X_10158_ _04488_ _04505_ _04507_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__and3_1
X_10089_ _04461_ _04463_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__xor2_1
X_13917_ clknet_leaf_72_clk _01136_ VGND VGND VPWR VPWR _122_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13848_ clknet_leaf_90_clk _01067_ VGND VGND VPWR VPWR _126_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13779_ clknet_leaf_94_clk _00998_ VGND VGND VPWR VPWR _130_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_clk clknet_3_2_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09941_ _03878_ _04320_ _01284_ _04321_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09872_ _04103_ _04110_ _03935_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__a21o_1
XFILLER_112_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _03179_ _03213_ _03212_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__o21ba_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08754_ _170_\[10\] _02801_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__and2_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07705_ _02208_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__inv_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08685_ _228_\[8\] _231_\[8\] VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_92_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _02160_ _02161_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__and2b_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07567_ _01675_ _01629_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__xnor2_1
X_06518_ _190_\[0\] _01215_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__or2_1
X_09306_ _185_\[27\] _03713_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__nand2_1
X_07498_ _02047_ _02048_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09237_ _03640_ _03642_ _03646_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__a21o_1
XFILLER_22_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09168_ _03578_ _03579_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__and2_1
X_09099_ _03493_ _03495_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__and2b_1
X_08119_ _234_\[11\] _02448_ _02636_ _02638_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__o211a_1
XFILLER_123_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11130_ _05226_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11061_ _164_\[25\] _04867_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__or2_1
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10012_ _04381_ _04389_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__nor2_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11963_ _05956_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_57_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13702_ clknet_leaf_59_clk _00921_ VGND VGND VPWR VPWR _134_\[6\] sky130_fd_sc_hd__dfxtp_1
X_11894_ _05897_ _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10914_ _164_\[6\] _167_\[6\] _05064_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__mux2_1
X_13633_ clknet_leaf_58_clk _00852_ VGND VGND VPWR VPWR _138_\[1\] sky130_fd_sc_hd__dfxtp_1
X_10845_ _170_\[18\] _05002_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__or2_1
XFILLER_13_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13564_ clknet_leaf_75_clk _00783_ VGND VGND VPWR VPWR _149_\[28\] sky130_fd_sc_hd__dfxtp_1
X_10776_ _170_\[30\] _173_\[30\] _04936_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__mux2_1
XFILLER_13_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13495_ clknet_leaf_41_clk _00714_ VGND VGND VPWR VPWR _158_\[13\] sky130_fd_sc_hd__dfxtp_1
X_12515_ _06294_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__clkbuf_1
X_12446_ _06200_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__buf_4
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12377_ _06222_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11328_ _152_\[19\] _05392_ _05318_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__mux2_1
XFILLER_5_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11259_ _05330_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__nand2_1
XFILLER_122_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_75_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08470_ _02889_ _02903_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__and2_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07421_ _01952_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__inv_2
XFILLER_51_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07352_ _01872_ _01893_ _01907_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__nand3_1
XFILLER_23_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07283_ _01839_ _01840_ _01838_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__a21o_1
XFILLER_31_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09022_ _01778_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__nor2_1
XFILLER_132_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09924_ _04210_ _04301_ _04302_ _04157_ _04305_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__o221a_1
XFILLER_120_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09855_ _04229_ _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__nor2_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08806_ _03218_ _03219_ _03227_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__or3b_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _04172_ _04173_ _03868_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__o21ai_1
X_06998_ _176_\[30\] _240_\[30\] _01569_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__mux2_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_16
X_08737_ _01974_ _03139_ _03161_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__o21a_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08668_ _02966_ _03092_ _03093_ _02965_ _03094_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__a2111o_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07619_ _02148_ _02165_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__nand2_1
XFILLER_54_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _173_\[18\] _176_\[18\] _01215_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__mux2_1
XFILLER_53_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08599_ _03027_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__xnor2_1
X_10561_ _173_\[27\] _04774_ _04835_ _04777_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__a211o_1
XFILLER_10_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12300_ _06181_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10492_ _176_\[7\] _04771_ _04751_ _04786_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__o211a_1
X_13280_ clknet_leaf_5_clk _00499_ VGND VGND VPWR VPWR _179_\[26\] sky130_fd_sc_hd__dfxtp_2
XFILLER_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12231_ _01393_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12162_ _140_\[9\] _138_\[9\] _06101_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__mux2_1
XFILLER_122_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12093_ _140_\[8\] _142_\[8\] _06068_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__mux2_1
X_11113_ _05213_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11044_ _164_\[18\] _01217_ _04627_ net45 _02833_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__o221a_1
XFILLER_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_16
X_12995_ clknet_leaf_15_clk _00214_ VGND VGND VPWR VPWR _240_\[3\] sky130_fd_sc_hd__dfxtp_1
X_11946_ _05944_ _05945_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__nand2_1
XFILLER_60_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11877_ _05883_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__clkbuf_1
X_13616_ clknet_leaf_47_clk _00835_ VGND VGND VPWR VPWR _140_\[16\] sky130_fd_sc_hd__dfxtp_2
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10828_ _167_\[13\] _04980_ _05009_ _05020_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__o211a_1
XFILLER_71_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13547_ clknet_leaf_84_clk _00766_ VGND VGND VPWR VPWR _149_\[11\] sky130_fd_sc_hd__dfxtp_1
X_10759_ _170_\[25\] _173_\[25\] _04936_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__mux2_1
XFILLER_145_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13478_ clknet_leaf_27_clk _00697_ _00111_ VGND VGND VPWR VPWR _190_\[0\] sky130_fd_sc_hd__dfrtp_1
X_12429_ _06249_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07970_ _01626_ _01608_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__xnor2_2
X_06921_ _240_\[7\] _01526_ _01510_ _01541_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__o211a_1
XFILLER_110_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09640_ _03901_ _03977_ _04032_ _03933_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__a211oi_1
X_06852_ _01448_ _01491_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__or2_1
XFILLER_95_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09571_ _03964_ _03966_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__xor2_1
X_06783_ _179_\[3\] _01299_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__or2_1
XFILLER_83_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_47_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_82_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08522_ _185_\[2\] _02913_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__nand2_1
XFILLER_91_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08453_ _02380_ _02883_ _02887_ _02202_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__o211a_1
XFILLER_36_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07404_ _01932_ _01933_ _01956_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__and3_1
XFILLER_51_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08384_ _02002_ _02831_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__or2_1
X_07335_ _01891_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__inv_2
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07266_ _01801_ _01819_ _01825_ _01799_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__o211a_1
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09005_ _03419_ _03421_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07197_ _01755_ _01758_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__xor2_1
XFILLER_3_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09907_ _04264_ _04265_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__or2_1
XFILLER_120_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09838_ _04222_ _04223_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__nand2_1
XFILLER_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09769_ _03910_ _01236_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__nand2_1
XFILLER_74_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _140_\[17\] _05812_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_38_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12780_ _122_\[15\] _120_\[15\] _06423_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__mux2_1
XFILLER_26_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _140_\[18\] _140_\[11\] VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__xnor2_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _05680_ _05683_ _05678_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__o21ai_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10613_ _173_\[11\] _04663_ _04871_ _04823_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__o211a_1
X_11593_ _118_\[21\] _118_\[25\] VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__xnor2_1
X_13401_ clknet_leaf_125_clk _00620_ VGND VGND VPWR VPWR _167_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13332_ clknet_leaf_9_clk _00551_ VGND VGND VPWR VPWR _173_\[14\] sky130_fd_sc_hd__dfxtp_1
X_10544_ _173_\[22\] _04818_ _04822_ _04823_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__o211a_1
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13263_ clknet_leaf_27_clk _00482_ VGND VGND VPWR VPWR _179_\[9\] sky130_fd_sc_hd__dfxtp_1
X_10475_ _04724_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__buf_2
XFILLER_6_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13194_ clknet_leaf_34_clk _00413_ VGND VGND VPWR VPWR _185_\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_142_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12214_ _06136_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12145_ _140_\[1\] _138_\[1\] _01394_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__mux2_1
X_12076_ _140_\[0\] _142_\[0\] _06005_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__mux2_1
XFILLER_96_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11027_ _03248_ _04861_ _05156_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__a21boi_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_29_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
X_12978_ clknet_leaf_23_clk _00197_ VGND VGND VPWR VPWR _243_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11929_ _142_\[18\] _05930_ _05893_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__mux2_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_28 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 _167_\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07120_ _237_\[26\] VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__buf_4
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07051_ _01615_ _01636_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__or2_1
XFILLER_127_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07953_ _02486_ _02487_ _02488_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__nand3_1
X_06904_ _01448_ _01529_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__or2_1
XFILLER_83_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07884_ _01707_ _02421_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__xnor2_4
X_09623_ _142_\[3\] _03974_ _04016_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__a21bo_1
X_06835_ _01444_ _01478_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__nand2_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09554_ _195_\[2\] _195_\[1\] VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__nand2_2
X_06766_ _01424_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09485_ _01277_ _03878_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__or2_1
XFILLER_64_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06697_ _01380_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__clkbuf_1
X_08505_ _02776_ _02937_ _01411_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__mux2_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08436_ net60 _01519_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__or2_1
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08367_ _02817_ _02791_ _02760_ _02818_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__o211a_1
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07318_ _01874_ _01875_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08298_ _164_\[31\] _228_\[31\] _02750_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__mux2_1
XFILLER_137_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07249_ _01807_ _01808_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__nand2_1
XFILLER_124_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10260_ _01212_ _04625_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__nand2_1
XFILLER_3_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10191_ _04437_ _03952_ _04026_ _04540_ _03894_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__o32a_1
XFILLER_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13950_ clknet_leaf_68_clk _01169_ VGND VGND VPWR VPWR _120_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12901_ clknet_leaf_90_clk _00125_ VGND VGND VPWR VPWR _116_\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13881_ clknet_leaf_90_clk _01100_ VGND VGND VPWR VPWR _124_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _118_\[8\] _120_\[8\] _06451_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__mux2_1
XFILLER_74_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _06424_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__clkbuf_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _05263_ _05735_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__nand2_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12694_ _124_\[6\] _122_\[6\] _06379_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__mux2_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11645_ _05672_ _05673_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 din[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlymetal6s2s_1
X_11576_ _05610_ _05611_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__nand2_1
Xinput15 din[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10527_ _173_\[17\] _04780_ _04811_ _04785_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__o211a_1
X_13315_ clknet_leaf_4_clk _00534_ VGND VGND VPWR VPWR _176_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13246_ clknet_leaf_7_clk _00465_ VGND VGND VPWR VPWR _182_\[24\] sky130_fd_sc_hd__dfxtp_1
X_10458_ _179_\[30\] _182_\[30\] _04743_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__mux2_1
XFILLER_6_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10389_ _179_\[10\] _182_\[10\] _04693_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__mux2_1
X_13177_ clknet_leaf_103_clk _00396_ VGND VGND VPWR VPWR _225_\[25\] sky130_fd_sc_hd__dfxtp_1
X_12128_ _06091_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__clkbuf_1
X_12059_ _152_\[30\] _06047_ _06048_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__nand3_1
XFILLER_84_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06620_ _01246_ _01306_ _01322_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__o21ba_1
XFILLER_92_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06551_ _158_\[12\] _01259_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__or2_1
XFILLER_92_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09270_ _03672_ _03674_ _03678_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__a21o_1
XFILLER_61_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08221_ _01417_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__buf_4
XFILLER_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08152_ _167_\[21\] _231_\[21\] _02626_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_9_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
X_08083_ _231_\[1\] _02611_ _01695_ _02612_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__o211a_1
X_07103_ _240_\[21\] _01660_ _01653_ _01677_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__o211a_1
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07034_ _173_\[6\] _01623_ _01617_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__mux2_1
XFILLER_134_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08985_ _170_\[17\] _02823_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__nand2_1
XFILLER_130_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07936_ _02471_ _02472_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__nand2_1
X_07867_ _182_\[24\] _01684_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__nand2_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09606_ _03998_ _03999_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__or2_1
X_06818_ _179_\[12\] _01299_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__or2_1
XFILLER_83_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07798_ _02308_ _02322_ _02338_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__o21ai_1
X_09537_ _01241_ _03896_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__nand2_1
X_06749_ _01408_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__buf_4
XFILLER_24_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09468_ _03866_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__inv_2
XFILLER_52_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09399_ _03762_ _03765_ _03803_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__a21oi_1
X_08419_ net55 _01519_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__or2_1
X_11430_ _116_\[1\] _05480_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11361_ _149_\[24\] _132_\[24\] VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10312_ _182_\[16\] _04634_ _04661_ _04649_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__o211a_1
XFILLER_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13100_ clknet_leaf_109_clk _00319_ VGND VGND VPWR VPWR _231_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11292_ _149_\[15\] _132_\[15\] VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__nand2_1
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10243_ _04605_ _04607_ _04604_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__a21oi_1
X_13031_ clknet_leaf_43_clk _00250_ VGND VGND VPWR VPWR _237_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10174_ _03899_ _04215_ _04544_ _03925_ _01233_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__o221a_1
XFILLER_3_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13933_ clknet_leaf_97_clk _01152_ VGND VGND VPWR VPWR _120_\[13\] sky130_fd_sc_hd__dfxtp_1
X_13864_ clknet_leaf_62_clk _01083_ VGND VGND VPWR VPWR _124_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12815_ _06004_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__clkbuf_4
X_13795_ clknet_leaf_63_clk _01014_ VGND VGND VPWR VPWR _128_\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _06415_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _01392_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__clkbuf_4
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11628_ _05646_ _05650_ _05658_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11559_ _05578_ _05580_ _05587_ _05596_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__o31a_1
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13229_ clknet_leaf_29_clk _00448_ VGND VGND VPWR VPWR _182_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08770_ _02037_ _03193_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__xnor2_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07721_ _185_\[20\] _234_\[20\] VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__nand2_1
X_07652_ _02164_ _02162_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__or2b_1
XFILLER_53_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06603_ _392_\[1\] _392_\[4\] _392_\[0\] VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__or3b_2
XFILLER_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07583_ _02129_ _02130_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__nor2_1
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06534_ _01242_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__buf_2
X_09322_ _03728_ _03729_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__and2b_1
XFILLER_34_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09253_ _170_\[25\] _02852_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__nand2_1
X_08204_ _164_\[4\] _02652_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__or2_1
X_09184_ _01923_ _03595_ _02002_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__a21o_1
X_08135_ _167_\[16\] _02616_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__or2_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08066_ _02595_ _02597_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__xnor2_4
XFILLER_108_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07017_ _01608_ _01565_ _01609_ _01610_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__o211a_1
XFILLER_115_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08968_ _185_\[16\] _03344_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__nand2_1
XFILLER_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08899_ _03316_ _03318_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__xor2_1
X_07919_ _02454_ _02455_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__nand2_1
XFILLER_84_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10930_ net37 _05068_ _05093_ _05086_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__a211o_1
XFILLER_29_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12600_ _128_\[25\] _126_\[25\] _06335_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__mux2_1
X_10861_ _167_\[22\] _05022_ _05043_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__o211a_1
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13580_ clknet_leaf_51_clk _00799_ VGND VGND VPWR VPWR _142_\[12\] sky130_fd_sc_hd__dfxtp_1
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10792_ _01213_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__buf_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ _130_\[24\] _128_\[24\] _06302_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__mux2_1
XFILLER_12_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12462_ _06266_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11413_ _149_\[29\] _132_\[29\] VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__nor2_1
X_12393_ _132_\[22\] _134_\[22\] _06230_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__mux2_1
X_11344_ _152_\[21\] _05406_ _05318_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__mux2_1
XFILLER_4_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11275_ _152_\[12\] _01368_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__and2_1
X_10226_ _03896_ _04132_ _03984_ _03878_ _01244_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__a32o_1
X_13014_ clknet_leaf_3_clk _00233_ VGND VGND VPWR VPWR _240_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10157_ _04527_ _04528_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__and2_1
XFILLER_94_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10088_ _142_\[23\] _04462_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13916_ clknet_leaf_72_clk _01135_ VGND VGND VPWR VPWR _122_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13847_ clknet_leaf_92_clk _01066_ VGND VGND VPWR VPWR _126_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13778_ clknet_leaf_94_clk _00997_ VGND VGND VPWR VPWR _130_\[18\] sky130_fd_sc_hd__dfxtp_1
X_12729_ _06406_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09940_ _01243_ _03904_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__nor2_1
X_09871_ _01231_ _01236_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__nand2_1
XFILLER_112_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _03243_ _03244_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__nand2_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08753_ _03172_ _03177_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__xor2_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07704_ _02246_ _02247_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__nand2_1
XFILLER_66_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08684_ _03109_ _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__xnor2_2
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07635_ _02179_ _02180_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__xnor2_4
XFILLER_80_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07566_ _02096_ _02097_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__and2b_1
XFILLER_41_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06517_ _190_\[1\] _01227_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__xnor2_1
X_09305_ _02865_ _03712_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07497_ _243_\[12\] _240_\[12\] _01642_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__mux2_2
X_09236_ _02422_ _03645_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__xor2_1
XFILLER_119_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09167_ _03573_ _03551_ _03577_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__nand3_1
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09098_ _03510_ _03511_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__xnor2_2
X_08118_ _02625_ _02637_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__or2_1
XFILLER_134_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08049_ _243_\[30\] _240_\[30\] _01704_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__mux2_4
XFILLER_122_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11060_ _03607_ _04855_ _04628_ net52 _05177_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__o221a_1
X_10011_ _04382_ _04384_ _04387_ _04388_ _04078_ _04210_ VGND VGND VPWR VPWR _04389_
+ sky130_fd_sc_hd__mux4_1
XFILLER_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13701_ clknet_leaf_59_clk _00920_ VGND VGND VPWR VPWR _134_\[5\] sky130_fd_sc_hd__dfxtp_1
X_11962_ _05959_ _05960_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__or2b_1
XFILLER_84_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11893_ _05888_ _05890_ _05886_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__o21ai_1
XFILLER_72_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10913_ net63 _05048_ _05081_ _05067_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__o211a_1
X_13632_ clknet_leaf_58_clk _00851_ VGND VGND VPWR VPWR _138_\[0\] sky130_fd_sc_hd__dfxtp_1
X_10844_ _164_\[17\] _05025_ _05032_ _05001_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__a211o_1
X_13563_ clknet_leaf_75_clk _00782_ VGND VGND VPWR VPWR _149_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10775_ _04671_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__clkbuf_4
X_12514_ _130_\[16\] _128_\[16\] _06291_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__mux2_1
X_13494_ clknet_leaf_41_clk _00713_ VGND VGND VPWR VPWR _158_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12445_ _06257_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12376_ _132_\[14\] _134_\[14\] _06219_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__mux2_1
XFILLER_60_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11327_ _05390_ _05391_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11258_ _05313_ _05323_ _05321_ _05320_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__a31o_1
XFILLER_95_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10209_ _04303_ _04103_ _04135_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__o21ai_1
X_11189_ _05271_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07420_ _01421_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__buf_4
XFILLER_62_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07351_ _01872_ _01893_ _01907_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07282_ _01838_ _01839_ _01840_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__nand3_1
XFILLER_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09021_ _03436_ _03437_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09923_ _01232_ _04280_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__or3b_1
XFILLER_140_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09854_ _04232_ _04234_ _04238_ _01237_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__o22a_1
XFILLER_112_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08805_ _03218_ _03219_ _03227_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__o21ba_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _04144_ _04151_ _04171_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__and3_1
XFILLER_100_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06997_ _243_\[29\] _01548_ _01545_ _01595_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__o211a_1
XFILLER_73_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _185_\[9\] _03138_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__nand2_1
XFILLER_39_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _02994_ _02995_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__nand2_1
XFILLER_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07618_ _02162_ _02164_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08598_ _02972_ _02976_ _02973_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__o21a_1
X_07549_ _02096_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10560_ _176_\[27\] _04833_ _04806_ _04834_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__o211a_1
XFILLER_10_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10491_ _179_\[7\] _04746_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__or2_1
X_09219_ _03562_ _03587_ _03629_ _03565_ _03588_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__o221a_1
X_12230_ _06144_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12161_ _06108_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12092_ _06072_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__clkbuf_1
X_11112_ _05212_ _158_\[5\] _05192_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__mux2_1
XFILLER_89_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11043_ net44 _04628_ _05167_ _05117_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__o211a_1
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_clk clknet_3_1_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12994_ clknet_leaf_15_clk _00213_ VGND VGND VPWR VPWR _240_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11945_ _152_\[20\] _05943_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__or2_1
XFILLER_91_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11876_ _142_\[13\] _05882_ _05765_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__mux2_1
X_13615_ clknet_leaf_45_clk _00834_ VGND VGND VPWR VPWR _140_\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10827_ _170_\[13\] _05002_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__or2_1
X_13546_ clknet_leaf_87_clk _00765_ VGND VGND VPWR VPWR _149_\[10\] sky130_fd_sc_hd__dfxtp_1
X_10758_ _04636_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__clkbuf_2
X_13477_ clknet_leaf_127_clk _00696_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfxtp_1
X_12428_ _132_\[7\] _130_\[7\] _06247_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__mux2_1
XFILLER_126_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10689_ _04685_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__buf_2
X_12359_ _132_\[6\] _134_\[6\] _06208_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__mux2_1
XFILLER_126_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06920_ _176_\[7\] _01531_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__or2_1
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06851_ _179_\[20\] _243_\[20\] _01449_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__mux2_1
X_09570_ _142_\[2\] _03965_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__xnor2_1
X_06782_ _01411_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__buf_4
XFILLER_95_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08521_ _02949_ _02952_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08452_ _02404_ _02886_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__nand2_1
XFILLER_36_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07403_ _01932_ _01933_ _01956_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__a21oi_1
X_08383_ net46 _02830_ _01353_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__mux2_1
X_07334_ _01889_ _01890_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07265_ _01409_ _01824_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__nand2_1
XFILLER_136_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09004_ _02192_ _03388_ _03420_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__a21oi_1
X_07196_ _01756_ _01757_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__nand2_1
XFILLER_144_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09906_ _04287_ _04288_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__or2b_1
XFILLER_101_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09837_ _04188_ _04191_ _04221_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__or3b_1
XFILLER_100_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _01243_ _03983_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__nor2_1
XFILLER_100_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08719_ _03105_ _03107_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__nor2_1
X_09699_ _04086_ _04089_ _03871_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__a21oi_1
X_11730_ _05749_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__clkbuf_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _116_\[25\] _05687_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__xnor2_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11592_ _05626_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__clkbuf_1
X_10612_ _02028_ _04870_ _04630_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__mux2_1
X_13400_ clknet_leaf_124_clk _00619_ VGND VGND VPWR VPWR _167_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13331_ clknet_leaf_23_clk _00550_ VGND VGND VPWR VPWR _173_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10543_ _01424_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13262_ clknet_leaf_26_clk _00481_ VGND VGND VPWR VPWR _179_\[8\] sky130_fd_sc_hd__dfxtp_1
X_10474_ _173_\[2\] _04725_ _04773_ _04728_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__a211o_1
X_13193_ clknet_leaf_34_clk _00412_ VGND VGND VPWR VPWR _185_\[3\] sky130_fd_sc_hd__dfxtp_2
X_12213_ _138_\[1\] _136_\[1\] _06134_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__mux2_1
X_12144_ _06099_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12075_ _142_\[31\] _05352_ _06062_ _06063_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__a22o_1
XFILLER_110_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11026_ _164_\[12\] _01217_ _04627_ net39 _02833_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__o221a_1
XFILLER_65_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12977_ clknet_leaf_14_clk _00196_ VGND VGND VPWR VPWR _243_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11928_ net10 _05929_ _05852_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__mux2_1
X_11859_ _152_\[12\] _05866_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__nand2_1
XFILLER_60_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_29 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 _170_\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13529_ clknet_leaf_47_clk _00748_ VGND VGND VPWR VPWR _152_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07050_ _173_\[10\] _01635_ _01617_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__mux2_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07952_ _185_\[27\] _234_\[27\] VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__nand2_1
X_06903_ _176_\[2\] _240_\[2\] _01449_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__mux2_1
XFILLER_68_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07883_ _01664_ _01616_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__xnor2_2
X_09622_ _03975_ _03987_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__or2b_1
X_06834_ _243_\[16\] _01438_ _01477_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__o21ai_1
XFILLER_83_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09553_ _01230_ _03932_ _03940_ _03922_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__o211a_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08504_ _02929_ _02930_ _02936_ _01269_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__a22o_1
X_06765_ _01423_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__buf_4
X_09484_ _03872_ _03881_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__nand2_1
XFILLER_102_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06696_ _118_\[13\] _116_\[13\] _01370_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__mux2_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08435_ _225_\[31\] VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__buf_4
XFILLER_24_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08366_ net42 _02798_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__or2_1
X_07317_ _243_\[6\] _240_\[6\] _01623_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__mux2_4
XFILLER_109_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08297_ _01480_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__clkbuf_4
XFILLER_125_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07248_ _185_\[4\] _234_\[4\] VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__or2_1
XFILLER_118_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07179_ _01736_ _01737_ _01269_ _01741_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10190_ _04558_ _04559_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__or2_1
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12900_ clknet_leaf_72_clk _00124_ VGND VGND VPWR VPWR _116_\[9\] sky130_fd_sc_hd__dfxtp_1
X_13880_ clknet_leaf_90_clk _01099_ VGND VGND VPWR VPWR _124_\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _06459_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__clkbuf_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _122_\[6\] _120_\[6\] _06423_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__mux2_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _06387_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__clkbuf_1
X_11713_ _05725_ _05731_ _05733_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__a21o_1
XFILLER_70_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _05665_ _05667_ _05663_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__o21ai_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 din[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
X_11575_ _116_\[16\] _05609_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__or2_1
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput16 din[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_10_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10526_ _04809_ _04810_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__or2_1
X_13314_ clknet_leaf_10_clk _00533_ VGND VGND VPWR VPWR _176_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13245_ clknet_leaf_5_clk _00464_ VGND VGND VPWR VPWR _182_\[23\] sky130_fd_sc_hd__dfxtp_2
X_10457_ _176_\[29\] _04735_ _04761_ _04740_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__o211a_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10388_ _04681_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__buf_2
XFILLER_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13176_ clknet_leaf_103_clk _00395_ VGND VGND VPWR VPWR _225_\[24\] sky130_fd_sc_hd__dfxtp_1
X_12127_ _140_\[24\] _142_\[24\] _06090_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__mux2_1
XFILLER_111_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12058_ _140_\[17\] _140_\[15\] VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__nand2_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11009_ net62 _04629_ _05146_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__o21a_1
XFILLER_65_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06550_ _158_\[11\] _158_\[10\] _01258_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__or3_1
XFILLER_80_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08220_ _231_\[8\] _02690_ _02664_ _02710_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__a211o_1
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08151_ _234_\[20\] _02659_ _02636_ _02661_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__o211a_1
XFILLER_134_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08082_ _167_\[1\] _01646_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__or2_1
X_07102_ _01670_ _01676_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__or2_1
X_07033_ _237_\[6\] VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__clkbuf_8
XFILLER_115_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08984_ _03398_ _03401_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07935_ _182_\[26\] _01690_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__nand2_1
XFILLER_29_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09605_ _142_\[4\] _03997_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__nor2_1
XFILLER_83_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07866_ _182_\[24\] _01684_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__or2_1
XFILLER_29_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06817_ _246_\[11\] _01407_ _01460_ _01465_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__a211o_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07797_ _02336_ _02337_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__xnor2_1
X_09536_ _01234_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__clkinv_2
X_06748_ _01269_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__buf_4
XFILLER_37_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09467_ _03866_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__inv_2
X_06679_ _01371_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__clkbuf_1
X_08418_ _225_\[27\] VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__buf_6
X_09398_ _03762_ _03765_ _03803_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__and3_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08349_ net38 _02798_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__or2_1
X_11360_ _05418_ _05420_ _152_\[23\] _05262_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_138_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10311_ _179_\[16\] _04646_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__or2_1
XFILLER_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13030_ clknet_leaf_42_clk _00249_ VGND VGND VPWR VPWR _237_\[6\] sky130_fd_sc_hd__dfxtp_1
X_11291_ _149_\[15\] _132_\[15\] VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__nor2_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10242_ _03946_ _04608_ _04609_ _00105_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__o211a_1
XFILLER_106_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10173_ _04437_ _04108_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__nand2_1
XFILLER_79_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13932_ clknet_leaf_97_clk _01151_ VGND VGND VPWR VPWR _120_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13863_ clknet_leaf_62_clk _01082_ VGND VGND VPWR VPWR _124_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13794_ clknet_leaf_63_clk _01013_ VGND VGND VPWR VPWR _128_\[2\] sky130_fd_sc_hd__dfxtp_1
X_12814_ _06450_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12745_ _124_\[30\] _122_\[30\] _06412_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__mux2_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12676_ _06378_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__clkbuf_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _05655_ _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__nand2_1
XFILLER_144_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11558_ _05576_ _05586_ _05585_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__a21o_1
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10509_ _173_\[12\] _04780_ _04798_ _04785_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__o211a_1
XFILLER_143_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11489_ _149_\[7\] _05532_ _05533_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__mux2_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13228_ clknet_leaf_28_clk _00447_ VGND VGND VPWR VPWR _182_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ clknet_leaf_111_clk _00378_ VGND VGND VPWR VPWR _225_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _185_\[20\] _234_\[20\] VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__or2_1
XFILLER_38_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07651_ _02195_ _02196_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__nor2_1
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06602_ _01302_ _01304_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__nor2_1
X_07582_ _02094_ _02114_ _02128_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__nor3_1
X_06533_ _01241_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__buf_2
XFILLER_80_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09321_ _03683_ _03707_ _03727_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09252_ _03659_ _03661_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__xor2_1
XFILLER_138_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09183_ _03593_ _03594_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__xor2_2
XFILLER_21_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08203_ _01437_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__clkbuf_4
XFILLER_119_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08134_ _01437_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__clkbuf_4
XFILLER_119_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08065_ _185_\[31\] _02596_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__xor2_4
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07016_ _173_\[2\] _01580_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__or2_1
XFILLER_142_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08967_ _02205_ _03384_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08898_ _02124_ _03280_ _03317_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__o21a_1
XFILLER_29_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07918_ _02452_ _02453_ _02451_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__a21o_1
XFILLER_90_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07849_ _02386_ _02387_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__nand2_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10860_ _170_\[22\] _05036_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__or2_1
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09519_ _03912_ _03916_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__xnor2_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10791_ _164_\[2\] _04983_ _04994_ _04939_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__o211a_1
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _06200_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__clkbuf_4
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12461_ _132_\[23\] _130_\[23\] _06258_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__mux2_1
XFILLER_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11412_ _05464_ _05465_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__or2b_1
XFILLER_40_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12392_ _06004_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__clkbuf_4
XFILLER_126_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11343_ _05404_ _05405_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11274_ _05343_ _05345_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__nand2_1
XFILLER_4_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10225_ _185_\[29\] _03870_ _03864_ _04593_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__o211a_1
X_13013_ clknet_leaf_3_clk _00232_ VGND VGND VPWR VPWR _240_\[21\] sky130_fd_sc_hd__dfxtp_1
X_10156_ _04495_ _04512_ _04526_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__or3_1
XFILLER_94_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10087_ _246_\[23\] _01316_ _04409_ _243_\[23\] _01499_ VGND VGND VPWR VPWR _04462_
+ sky130_fd_sc_hd__o221a_1
XFILLER_47_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13915_ clknet_leaf_90_clk _01134_ VGND VGND VPWR VPWR _122_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13846_ clknet_leaf_92_clk _01065_ VGND VGND VPWR VPWR _126_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10989_ net56 _05110_ _05134_ _05122_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__a211o_1
XFILLER_15_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13777_ clknet_leaf_95_clk _00996_ VGND VGND VPWR VPWR _130_\[17\] sky130_fd_sc_hd__dfxtp_1
X_12728_ _124_\[22\] _122_\[22\] _06401_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__mux2_1
X_12659_ _126_\[21\] _124_\[21\] _06368_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__mux2_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09870_ _01243_ _04010_ _03936_ _04253_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__o31a_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _170_\[12\] _02807_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__nand2_1
XFILLER_85_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _03100_ _03173_ _03176_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__o21ai_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08683_ _01904_ _01905_ _03077_ _03076_ _03074_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__o32a_2
XFILLER_66_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07703_ _02242_ _02245_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__nand2_1
X_07634_ _02169_ _02173_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__or2_2
XFILLER_54_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07565_ _01650_ _01827_ _01693_ _02113_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__a211o_1
XFILLER_22_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06516_ _190_\[0\] _01226_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__nand2_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07496_ _02045_ _02046_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__or2_1
X_09304_ _02823_ _02794_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09235_ _185_\[25\] _03644_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09166_ _03573_ _03551_ _03577_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__a21o_1
XFILLER_134_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09097_ _170_\[20\] _02835_ _03476_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__a21o_1
X_08117_ _167_\[11\] _231_\[11\] _02626_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__mux2_1
XFILLER_123_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08048_ _02579_ _02580_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__or2b_1
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10010_ _03876_ _03893_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__nor2_1
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09999_ _243_\[20\] _04129_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__or2_1
XFILLER_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11961_ _152_\[21\] _05958_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__nand2_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13700_ clknet_leaf_58_clk _00919_ VGND VGND VPWR VPWR _134_\[4\] sky130_fd_sc_hd__dfxtp_1
X_10912_ _05079_ _05080_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__or2_1
XFILLER_17_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11892_ _152_\[15\] _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13631_ clknet_leaf_53_clk _00850_ VGND VGND VPWR VPWR _140_\[31\] sky130_fd_sc_hd__dfxtp_2
X_10843_ _167_\[17\] _05022_ _05009_ _05031_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__o211a_1
X_13562_ clknet_leaf_75_clk _00781_ VGND VGND VPWR VPWR _149_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10774_ _167_\[29\] _04945_ _04982_ _04952_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__a211o_1
XFILLER_12_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12513_ _06293_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__clkbuf_1
X_13493_ clknet_leaf_46_clk _00712_ VGND VGND VPWR VPWR _158_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12444_ _132_\[15\] _130_\[15\] _06247_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__mux2_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12375_ _06221_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11326_ _05381_ _05386_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__nand2_1
XFILLER_4_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11257_ _05313_ _05323_ _05321_ _05330_ _05320_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__a311o_2
XFILLER_106_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10208_ _04303_ _04085_ _04576_ _01239_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__o211a_1
X_11188_ _152_\[1\] _05270_ _01362_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__mux2_1
X_10139_ _03946_ _04510_ _04511_ _00105_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__o211a_1
XFILLER_79_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13829_ clknet_leaf_63_clk _01048_ VGND VGND VPWR VPWR _126_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07350_ _01903_ _01906_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__xor2_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07281_ _185_\[5\] _234_\[5\] VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__nand2_1
X_09020_ _03404_ _03406_ _03403_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__a21bo_1
XFILLER_116_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09922_ _04075_ _01285_ _03875_ _04303_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__or4_1
X_09853_ _03871_ _03897_ _04235_ _04237_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__o31a_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _04144_ _04151_ _04171_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__a21oi_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08804_ _02048_ _03226_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _01568_ _01594_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__or2_1
X_08735_ _02006_ _03159_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__xnor2_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _03020_ _03021_ _03050_ _03086_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__nand4b_1
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _02123_ _02125_ _02163_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__o21ba_1
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08597_ _03025_ _03026_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__nand2_1
XFILLER_14_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07548_ _243_\[14\] _240_\[14\] _01650_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__mux2_2
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07479_ _01638_ _01973_ _01886_ _02030_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__o211a_1
XFILLER_22_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10490_ _173_\[6\] _04780_ _04784_ _04785_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__o211a_1
X_09218_ _03564_ _03589_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__nand2_1
XFILLER_10_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09149_ _03545_ _03546_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__o21ai_1
X_12160_ _140_\[8\] _138_\[8\] _06101_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__mux2_1
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11111_ net6 _05211_ _05196_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__mux2_1
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12091_ _140_\[7\] _142_\[7\] _06068_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__mux2_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11042_ _164_\[17\] _04865_ _04638_ _05166_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__a211o_1
XFILLER_131_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12993_ clknet_leaf_17_clk _00212_ VGND VGND VPWR VPWR _240_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11944_ _152_\[20\] _05943_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__nand2_1
XFILLER_45_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11875_ net5 _05881_ _05852_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__mux2_1
XFILLER_72_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13614_ clknet_leaf_49_clk _00833_ VGND VGND VPWR VPWR _140_\[14\] sky130_fd_sc_hd__dfxtp_2
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10826_ _164_\[12\] _04986_ _05019_ _05001_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__a211o_1
XFILLER_111_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13545_ clknet_leaf_68_clk _00764_ VGND VGND VPWR VPWR _149_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10757_ _167_\[24\] _04945_ _04970_ _04952_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__a211o_1
XFILLER_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10688_ _167_\[4\] _04836_ _04921_ _04914_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__a211o_1
XFILLER_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13476_ clknet_leaf_126_clk _00695_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_1
X_12427_ _06248_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12358_ _06212_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12289_ _06175_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11309_ _149_\[17\] _132_\[17\] VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__nand2_1
XFILLER_141_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06850_ _246_\[19\] _01485_ _01481_ _01490_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__o211a_1
XFILLER_95_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06781_ _01437_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__clkbuf_4
XFILLER_82_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08520_ _185_\[3\] _02951_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08451_ _02884_ _02885_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__nand2_1
XFILLER_36_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07402_ _01952_ _01955_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__xor2_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08382_ _225_\[19\] VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__buf_4
XFILLER_32_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07333_ _01859_ _01862_ _01858_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__o21a_1
XFILLER_50_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_124_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_124_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07264_ _01822_ _01823_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__xnor2_2
XFILLER_31_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09003_ _03385_ _03387_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__nor2_1
XFILLER_117_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07195_ _185_\[2\] _234_\[2\] VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__or2_1
XFILLER_144_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09905_ _04250_ _04262_ _04286_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__o21ai_1
XFILLER_101_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09836_ _04188_ _04191_ _04221_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__o21bai_2
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _04153_ _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__or2_1
XFILLER_100_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06979_ _01495_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__buf_2
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09698_ _03983_ _04087_ _04088_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__a21oi_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _01960_ _03143_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__xnor2_2
XFILLER_27_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _03074_ _03076_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__xnor2_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _118_\[11\] _05686_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__xnor2_2
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11591_ _149_\[17\] _05624_ _05625_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__mux2_1
X_10611_ _176_\[11\] _04867_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__or2_1
XFILLER_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_115_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_115_clk sky130_fd_sc_hd__clkbuf_16
X_13330_ clknet_leaf_23_clk _00549_ VGND VGND VPWR VPWR _173_\[12\] sky130_fd_sc_hd__dfxtp_1
X_10542_ _04809_ _04821_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__or2_1
X_13261_ clknet_leaf_29_clk _00480_ VGND VGND VPWR VPWR _179_\[7\] sky130_fd_sc_hd__dfxtp_1
X_12212_ _06135_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10473_ _176_\[2\] _04771_ _04751_ _04772_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__o211a_1
X_13192_ clknet_leaf_34_clk _00411_ VGND VGND VPWR VPWR _185_\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_108_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12143_ _140_\[0\] _138_\[0\] _01394_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__mux2_1
XFILLER_123_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12074_ net25 _05742_ _05263_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__o21a_1
XFILLER_97_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11025_ net38 _04628_ _05155_ _05117_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__o211a_1
XFILLER_77_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12976_ clknet_leaf_14_clk _00195_ VGND VGND VPWR VPWR _243_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11927_ _05924_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__xor2_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11858_ _140_\[22\] _05865_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11789_ _140_\[23\] _05802_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__xnor2_1
XANTENNA_19 _170_\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10809_ _04971_ _05007_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_106_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_106_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13528_ clknet_leaf_47_clk _00747_ VGND VGND VPWR VPWR _152_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13459_ clknet_leaf_123_clk _00678_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_2
XFILLER_133_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_776 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07951_ _185_\[27\] _234_\[27\] VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__or2_1
X_06902_ _243_\[1\] _01496_ _01509_ _01528_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__a211o_1
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07882_ _02391_ _02392_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__and2b_1
X_09621_ _04000_ _04014_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__xnor2_1
X_06833_ _179_\[16\] _01301_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__or2_1
XFILLER_68_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09552_ _142_\[1\] _03921_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__and2_1
X_06764_ _01416_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__inv_2
XFILLER_102_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08503_ _02932_ _02935_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__xnor2_1
X_09483_ _03873_ _03876_ _03878_ _03880_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__a22o_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06695_ _01379_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08434_ _228_\[30\] _02845_ _02834_ _02870_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__o211a_1
XFILLER_24_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08365_ _225_\[15\] VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__buf_4
X_07316_ _01872_ _01873_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__nand2_1
XFILLER_137_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08296_ _231_\[30\] _02706_ _02695_ _02764_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__o211a_1
X_07247_ _185_\[4\] _234_\[4\] VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_2_0_clk clknet_3_1_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_117_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07178_ _01711_ _01740_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09819_ _04195_ _04202_ _04204_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__and3_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12830_ _118_\[7\] _120_\[7\] _06451_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__mux2_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _01392_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__clkbuf_8
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12692_ _124_\[5\] _122_\[5\] _06379_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__mux2_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _05725_ _05731_ _05733_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__and3_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11643_ _116_\[23\] _05671_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__xnor2_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput17 din[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
Xinput28 din[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
X_11574_ _116_\[16\] _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__nand2_1
XFILLER_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10525_ _176_\[17\] _179_\[17\] _04790_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__mux2_1
X_13313_ clknet_leaf_8_clk _00532_ VGND VGND VPWR VPWR _176_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13244_ clknet_leaf_6_clk _00463_ VGND VGND VPWR VPWR _182_\[22\] sky130_fd_sc_hd__dfxtp_1
X_10456_ _04712_ _04760_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__or2_1
XFILLER_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13175_ clknet_leaf_101_clk _00394_ VGND VGND VPWR VPWR _225_\[23\] sky130_fd_sc_hd__dfxtp_1
X_12126_ _06004_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__buf_4
X_10387_ _176_\[9\] _04691_ _04711_ _04677_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__o211a_1
XFILLER_111_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12057_ _140_\[17\] _140_\[15\] VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__or2_1
XFILLER_77_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11008_ _164_\[4\] _04678_ _02977_ _04686_ _04648_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__o221a_1
XFILLER_38_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12959_ clknet_leaf_20_clk _00178_ VGND VGND VPWR VPWR _246_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08150_ _02625_ _02660_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__or2_1
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07101_ _173_\[21\] _01675_ _01672_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__mux2_1
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08081_ _01437_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__clkbuf_4
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07032_ _240_\[5\] _01601_ _01598_ _01622_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__o211a_1
XFILLER_127_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08983_ _03399_ _03368_ _03400_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__o21ai_1
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07934_ _182_\[26\] _01690_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__or2_1
XFILLER_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07865_ _01408_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__clkbuf_4
XFILLER_29_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09604_ _142_\[4\] _03997_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__and2_1
XFILLER_110_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06816_ _243_\[11\] _01438_ _01461_ _01464_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__o211a_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07796_ _243_\[22\] _240_\[22\] _01678_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__mux2_4
X_09535_ _01234_ _03898_ _03926_ _03931_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__a31o_1
X_06747_ _01406_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__clkbuf_4
XFILLER_71_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09466_ _03866_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__inv_2
X_06678_ _118_\[4\] _116_\[4\] _01370_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__mux2_1
XFILLER_52_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08417_ _228_\[26\] _02845_ _02834_ _02857_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__o211a_1
XFILLER_24_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09397_ _03801_ _03802_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__nor2_1
XFILLER_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08348_ _225_\[11\] VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__clkbuf_4
X_08279_ _231_\[25\] _02706_ _02695_ _02752_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__o211a_1
XFILLER_125_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11290_ _05359_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__clkbuf_1
X_10310_ _179_\[15\] _04658_ _04660_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__a21o_1
X_10241_ _185_\[30\] _03867_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__or2_1
XFILLER_4_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10172_ _03954_ _04156_ _04542_ _01238_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__a211o_1
XFILLER_121_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13931_ clknet_leaf_96_clk _01150_ VGND VGND VPWR VPWR _120_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13862_ clknet_leaf_62_clk _01081_ VGND VGND VPWR VPWR _124_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13793_ clknet_leaf_63_clk _01012_ VGND VGND VPWR VPWR _128_\[1\] sky130_fd_sc_hd__dfxtp_1
X_12813_ _122_\[31\] _120_\[31\] _01367_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__mux2_1
XFILLER_62_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12744_ _06414_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__clkbuf_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12675_ _126_\[29\] _124_\[29\] _06368_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__mux2_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11626_ _05656_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__inv_2
X_11557_ _05593_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__nand2_1
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10508_ _04766_ _04797_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__or2_1
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11488_ _01361_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__buf_4
XFILLER_6_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13227_ clknet_leaf_29_clk _00446_ VGND VGND VPWR VPWR _182_\[5\] sky130_fd_sc_hd__dfxtp_1
X_10439_ _182_\[24\] _04746_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__or2_1
XFILLER_124_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ clknet_leaf_109_clk _00377_ VGND VGND VPWR VPWR _225_\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12109_ _06081_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13089_ clknet_leaf_111_clk _00308_ VGND VGND VPWR VPWR _231_\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07650_ _02158_ _02182_ _02193_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__nor3_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06601_ _01303_ _01297_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__nor2_1
XFILLER_92_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07581_ _02094_ _02114_ _02128_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__o21a_1
X_06532_ _01240_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__clkbuf_4
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09320_ _03683_ _03707_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__nor3_1
X_09251_ _03628_ _03634_ _03660_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__a21bo_1
XFILLER_61_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08202_ _231_\[3\] _02659_ _02695_ _02697_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__o211a_1
XFILLER_119_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09182_ _03541_ _03543_ _03540_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__a21o_1
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08133_ _234_\[15\] _02646_ _02629_ _02648_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__a211o_1
XFILLER_119_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08064_ _243_\[31\] _240_\[31\] _01707_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__mux2_2
X_07015_ _01420_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__buf_2
XFILLER_108_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08966_ _185_\[17\] _03383_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08897_ _185_\[14\] _03279_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__nand2_1
X_07917_ _02451_ _02452_ _02453_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_95_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07848_ _02384_ _02385_ _02383_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__a21o_1
X_09518_ _142_\[0\] _03915_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__xnor2_1
X_07779_ _01856_ _02300_ _02320_ _01884_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__a211o_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10790_ _04971_ _04993_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__or2_1
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09449_ _02839_ _03852_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12460_ _06265_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11411_ _149_\[30\] _132_\[30\] VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__or2_1
X_12391_ _06229_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11342_ _05395_ _05400_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__nand2_1
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11273_ _05328_ _05331_ _05336_ _05335_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__a31o_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10224_ _03945_ _04591_ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__or3_1
XFILLER_106_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13012_ clknet_leaf_3_clk _00231_ VGND VGND VPWR VPWR _240_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10155_ _04495_ _04512_ _04526_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__o21ai_1
XFILLER_79_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10086_ _04054_ _04456_ _04457_ _04460_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_86_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_16
X_13914_ clknet_leaf_91_clk _01133_ VGND VGND VPWR VPWR _122_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13845_ clknet_leaf_93_clk _01064_ VGND VGND VPWR VPWR _126_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13776_ clknet_leaf_93_clk _00995_ VGND VGND VPWR VPWR _130_\[16\] sky130_fd_sc_hd__dfxtp_1
X_10988_ _164_\[28\] _05107_ _04865_ _05133_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__o211a_1
X_12727_ _06405_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12658_ _06369_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__clkbuf_1
X_11609_ _05629_ _05634_ _05641_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_10_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
X_12589_ _128_\[20\] _126_\[20\] _06324_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__mux2_1
XFILLER_144_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _170_\[12\] _02807_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__or2_1
XFILLER_98_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08751_ _03134_ _03174_ _03175_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__a21o_1
XFILLER_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08682_ _01939_ _03108_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__xnor2_4
XFILLER_66_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07702_ _02242_ _02245_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__or2_1
XFILLER_93_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07633_ _182_\[17\] _01661_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__xnor2_2
XFILLER_53_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07564_ _01801_ _02105_ _02112_ _01799_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__o211a_1
XFILLER_41_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07495_ _02011_ _02038_ _02044_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__and3_1
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09303_ _02451_ _03710_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__nand2_1
XFILLER_22_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06515_ _01225_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__buf_6
X_09234_ _02858_ _03643_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09165_ _02362_ _03576_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__xor2_1
XFILLER_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08116_ _01480_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__clkbuf_4
XFILLER_135_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09096_ _03508_ _03509_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__nand2_1
XFILLER_116_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08047_ _02578_ _02577_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09998_ _04358_ _04369_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__nor2_1
XFILLER_76_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08949_ _03367_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_68_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_16
X_11960_ _152_\[21\] _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__nor2_1
XFILLER_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10911_ _164_\[5\] _167_\[5\] _05064_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__mux2_1
XFILLER_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11891_ _140_\[25\] _05895_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__xnor2_2
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13630_ clknet_leaf_51_clk _00849_ VGND VGND VPWR VPWR _140_\[30\] sky130_fd_sc_hd__dfxtp_2
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10842_ _170_\[17\] _05002_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__or2_1
X_13561_ clknet_leaf_75_clk _00780_ VGND VGND VPWR VPWR _149_\[25\] sky130_fd_sc_hd__dfxtp_1
X_10773_ _170_\[29\] _04980_ _04958_ _04981_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__o211a_1
XFILLER_25_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12512_ _130_\[15\] _128_\[15\] _06291_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__mux2_1
X_13492_ clknet_leaf_46_clk _00711_ VGND VGND VPWR VPWR _158_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12443_ _06256_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__clkbuf_1
X_12374_ _132_\[13\] _134_\[13\] _06219_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__mux2_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11325_ _05388_ _05389_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__or2b_1
X_11256_ _05329_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__inv_2
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10207_ _03890_ _03927_ _01244_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__a21o_1
X_11187_ _05264_ _05269_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10138_ _185_\[25\] _03867_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__or2_1
XFILLER_95_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_59_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_16
X_10069_ _04434_ _04443_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__nand2_1
XFILLER_48_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13828_ clknet_leaf_63_clk _01047_ VGND VGND VPWR VPWR _126_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13759_ clknet_leaf_57_clk _00978_ VGND VGND VPWR VPWR _132_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07280_ _185_\[5\] _234_\[5\] VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__or2_1
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09921_ _01278_ _01281_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__nor2_2
XFILLER_104_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09852_ _03910_ _03906_ _04236_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__or3_1
XFILLER_112_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09783_ _04169_ _04170_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08803_ _03223_ _03225_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__xor2_1
XFILLER_58_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _185_\[10\] _03158_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__xnor2_1
X_06995_ _176_\[29\] _240_\[29\] _01569_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__mux2_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _02904_ _02928_ _02964_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07616_ _02126_ _02127_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__and2b_1
X_08596_ _170_\[5\] _02784_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__nand2_1
X_07547_ _02094_ _02095_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__or2_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07478_ _02022_ _02023_ _02029_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__o21ai_1
XFILLER_22_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09217_ _03625_ _03627_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09148_ _03558_ _03560_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__xnor2_1
X_09079_ _228_\[20\] _231_\[20\] _02835_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__a21o_1
X_11110_ _01255_ _05210_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__nand2_1
XFILLER_107_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12090_ _06071_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11041_ _03407_ _04630_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__nor2_1
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12992_ clknet_leaf_17_clk _00211_ VGND VGND VPWR VPWR _240_\[0\] sky130_fd_sc_hd__dfxtp_1
X_11943_ _140_\[30\] _05942_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11874_ _05879_ _05880_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__xnor2_1
X_13613_ clknet_leaf_51_clk _00832_ VGND VGND VPWR VPWR _140_\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_44_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10825_ _167_\[12\] _04980_ _05009_ _05018_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__o211a_1
XFILLER_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13544_ clknet_leaf_74_clk _00763_ VGND VGND VPWR VPWR _149_\[8\] sky130_fd_sc_hd__dfxtp_1
X_10756_ _170_\[24\] _04942_ _04958_ _04969_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__o211a_1
XFILLER_139_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10687_ _170_\[4\] _04833_ _04806_ _04920_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__o211a_1
XFILLER_9_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13475_ clknet_leaf_122_clk _00694_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_2
XFILLER_139_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12426_ _132_\[6\] _130_\[6\] _06247_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__mux2_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12357_ _132_\[5\] _134_\[5\] _06208_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__mux2_1
X_12288_ _136_\[5\] _134_\[5\] _06167_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__mux2_1
XFILLER_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11308_ _149_\[17\] _132_\[17\] VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__nor2_1
XFILLER_141_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11239_ _149_\[6\] _132_\[6\] _05306_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__nand3_1
XFILLER_110_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06780_ _01408_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__buf_4
XFILLER_82_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08450_ _170_\[0\] _02768_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__or2_1
XFILLER_36_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07401_ _01953_ _01954_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__nand2_1
X_08381_ _228_\[18\] _02775_ _02810_ _02829_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__a211o_1
X_07332_ _01887_ _01888_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__nand2_1
XFILLER_16_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07263_ _01749_ _01772_ _01775_ _01773_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__o31a_2
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07194_ _185_\[2\] _234_\[2\] VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__nand2_1
X_09002_ _02216_ _03418_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09904_ _04250_ _04262_ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__nor3_1
XFILLER_104_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09835_ _04219_ _04220_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__or2_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _142_\[10\] _04152_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__nor2_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06978_ _243_\[23\] _01536_ _01557_ _01582_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__a211o_1
XFILLER_46_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09697_ _01234_ _03884_ _03903_ _03928_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__and4_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08717_ _03140_ _03142_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__xnor2_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _03033_ _03036_ _03075_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__o21a_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _185_\[4\] _02981_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__nand2_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11590_ _01361_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__buf_4
X_10610_ _173_\[10\] _04663_ _04869_ _04823_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__o211a_1
XFILLER_50_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10541_ _176_\[22\] _179_\[22\] _04790_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__mux2_1
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13260_ clknet_leaf_28_clk _00479_ VGND VGND VPWR VPWR _179_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12211_ _138_\[0\] _136_\[0\] _06134_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__mux2_1
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10472_ _179_\[2\] _04746_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__or2_1
XFILLER_41_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13191_ clknet_leaf_34_clk _00410_ VGND VGND VPWR VPWR _185_\[1\] sky130_fd_sc_hd__dfxtp_2
X_12142_ _06098_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12073_ _06049_ _06055_ _06060_ _06061_ _05776_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__a311o_1
XFILLER_110_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11024_ _164_\[11\] _04865_ _04638_ _05154_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__a211o_1
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12975_ clknet_leaf_18_clk _00194_ VGND VGND VPWR VPWR _243_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11926_ _05909_ _05925_ _05927_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__o21a_1
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11857_ _140_\[29\] _140_\[31\] VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11788_ _140_\[25\] _140_\[16\] VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10808_ _167_\[7\] _170_\[7\] _04995_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__mux2_1
X_13527_ clknet_leaf_76_clk _00746_ VGND VGND VPWR VPWR _152_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10739_ _04685_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__clkbuf_4
XFILLER_118_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13458_ clknet_leaf_114_clk _00677_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_2
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12409_ _132_\[30\] _134_\[30\] _06230_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__mux2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13389_ clknet_leaf_1_clk _00608_ VGND VGND VPWR VPWR _167_\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_127_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07950_ _01671_ _02485_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__xnor2_4
XFILLER_141_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06901_ _240_\[1\] _01526_ _01510_ _01527_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__o211a_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07881_ _01480_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__clkbuf_4
X_09620_ _04008_ _04013_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__or2_1
X_06832_ _246_\[15\] _01407_ _01460_ _01476_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__a211o_1
XFILLER_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09551_ _185_\[1\] _03869_ _03919_ _03947_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__o211a_1
XFILLER_110_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06763_ _01421_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__buf_2
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08502_ _02933_ _02934_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__nor2_1
X_09482_ _03879_ _03875_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__nor2_4
XFILLER_91_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06694_ _118_\[12\] _116_\[12\] _01370_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__mux2_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08433_ _02002_ _02869_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__or2_1
XFILLER_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08364_ _228_\[14\] _02771_ _02765_ _02816_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__o211a_1
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07315_ _01840_ _01841_ _01871_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__nand3_1
XFILLER_32_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08295_ _02749_ _02763_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__or2_1
X_07246_ _01701_ _01805_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__xnor2_1
X_07177_ _01738_ _01739_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__nor2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09818_ _04197_ _04194_ _04201_ _04203_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_101_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09749_ _01284_ _03903_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__nor2_1
XFILLER_101_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _06422_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__clkbuf_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12691_ _06386_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__clkbuf_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _116_\[30\] _05732_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__xor2_1
XFILLER_70_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11642_ _118_\[9\] _05670_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__xnor2_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput18 din[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
X_11573_ _118_\[19\] _05608_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__xnor2_1
X_13312_ clknet_leaf_5_clk _00531_ VGND VGND VPWR VPWR _176_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput29 din[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10524_ _04681_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__buf_2
XFILLER_136_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13243_ clknet_leaf_6_clk _00462_ VGND VGND VPWR VPWR _182_\[21\] sky130_fd_sc_hd__dfxtp_1
X_10455_ _179_\[29\] _182_\[29\] _04743_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__mux2_1
X_13174_ clknet_leaf_103_clk _00393_ VGND VGND VPWR VPWR _225_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12125_ _06089_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__clkbuf_1
X_10386_ _04692_ _04710_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__or2_1
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12056_ _06046_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11007_ net61 _04629_ _05145_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__o21a_1
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12958_ clknet_leaf_22_clk _00177_ VGND VGND VPWR VPWR _246_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12889_ _04648_ _06490_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__and2_1
X_11909_ _05912_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07100_ _237_\[21\] VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__buf_6
X_08080_ _234_\[0\] _02448_ _02419_ _02610_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__o211a_1
X_07031_ _01615_ _01621_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__or2_1
XFILLER_127_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08982_ _03358_ _03357_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__or2b_1
XFILLER_114_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07933_ _02467_ _02468_ _02465_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__o21ai_1
XFILLER_96_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07864_ _02396_ _02402_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__xnor2_1
XFILLER_113_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09603_ _246_\[4\] _01313_ _03913_ _243_\[4\] _01442_ VGND VGND VPWR VPWR _03997_
+ sky130_fd_sc_hd__o221a_1
X_06815_ _179_\[11\] _01299_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__or2_1
XFILLER_68_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07795_ _02334_ _02335_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__or2_1
X_09534_ _01241_ _03903_ _03927_ _03930_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__a31oi_1
X_06746_ _01405_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__buf_4
XFILLER_64_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09465_ _03866_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__inv_2
X_06677_ _01367_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__buf_4
X_08416_ _02002_ _02856_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__or2_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09396_ _03756_ _03777_ _03799_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__nor3_1
XFILLER_12_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08347_ _228_\[10\] _02775_ _02753_ _02803_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__a211o_1
X_08278_ _02749_ _02751_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__or2_1
XFILLER_137_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07229_ _01788_ _01789_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10240_ _04606_ _04607_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__xor2_1
XFILLER_106_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10171_ _04081_ _04010_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__nor2_1
XFILLER_121_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13930_ clknet_leaf_97_clk _01149_ VGND VGND VPWR VPWR _120_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13861_ clknet_leaf_64_clk _01080_ VGND VGND VPWR VPWR _124_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13792_ clknet_leaf_65_clk _01011_ VGND VGND VPWR VPWR _128_\[0\] sky130_fd_sc_hd__dfxtp_1
X_12812_ _06449_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12743_ _124_\[29\] _122_\[29\] _06412_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__mux2_1
XFILLER_55_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12674_ _06377_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__clkbuf_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11625_ _116_\[21\] _05654_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__nor2_1
X_11556_ _116_\[14\] _05592_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__or2_1
XFILLER_11_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10507_ _176_\[12\] _179_\[12\] _04790_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__mux2_1
X_13226_ clknet_leaf_27_clk _00445_ VGND VGND VPWR VPWR _182_\[4\] sky130_fd_sc_hd__dfxtp_1
X_11487_ _05530_ _05531_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10438_ _176_\[23\] _04725_ _04748_ _04728_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__a211o_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10369_ _179_\[4\] _182_\[4\] _04693_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__mux2_1
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ clknet_leaf_111_clk _00376_ VGND VGND VPWR VPWR _225_\[5\] sky130_fd_sc_hd__dfxtp_1
X_12108_ _140_\[15\] _142_\[15\] _06079_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__mux2_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13088_ clknet_leaf_115_clk _00307_ VGND VGND VPWR VPWR _231_\[0\] sky130_fd_sc_hd__dfxtp_1
X_12039_ _140_\[13\] _140_\[15\] VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__xor2_1
XFILLER_78_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_1_0_clk clknet_3_0_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_06600_ net35 VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__inv_2
XFILLER_93_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07580_ _02126_ _02127_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__xnor2_1
X_06531_ _195_\[3\] VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__buf_2
XFILLER_81_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09250_ _03627_ _03625_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__or2b_1
XFILLER_21_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08201_ _02686_ _02696_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__or2_1
X_09181_ _170_\[23\] _02846_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__xor2_2
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08132_ _231_\[15\] _02611_ _02641_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__o211a_1
X_08063_ _01684_ _02594_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__xnor2_2
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07014_ _237_\[2\] VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__buf_4
XFILLER_134_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08965_ _02868_ _03382_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07916_ _185_\[26\] _234_\[26\] VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__nand2_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08896_ _02117_ _03315_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07847_ _02383_ _02384_ _02385_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__nand3_1
XFILLER_83_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07778_ _02316_ _02318_ _02319_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__o21a_1
XFILLER_44_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09517_ _246_\[0\] _01314_ _03914_ _243_\[0\] _01413_ VGND VGND VPWR VPWR _03915_
+ sky130_fd_sc_hd__o221a_2
X_06729_ _01398_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _03814_ _03819_ _03817_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__o21ai_1
XFILLER_138_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09379_ _02540_ _03784_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__nand2_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11410_ _149_\[30\] _132_\[30\] VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__and2_1
X_12390_ _132_\[21\] _134_\[21\] _06219_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__mux2_1
XFILLER_126_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11341_ _05402_ _05403_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__or2b_1
XFILLER_141_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11272_ _05328_ _05331_ _05336_ _05343_ _05335_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__a311o_2
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10223_ _04572_ _04568_ _04590_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__o21a_1
X_13011_ clknet_leaf_9_clk _00230_ VGND VGND VPWR VPWR _240_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10154_ _04524_ _04525_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10085_ _01238_ _04458_ _04459_ _01232_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__o211a_1
XFILLER_87_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13913_ clknet_leaf_91_clk _01132_ VGND VGND VPWR VPWR _122_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13844_ clknet_leaf_93_clk _01063_ VGND VGND VPWR VPWR _126_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13775_ clknet_leaf_84_clk _00994_ VGND VGND VPWR VPWR _130_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10987_ _167_\[28\] _04867_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__or2_1
XFILLER_16_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12726_ _124_\[21\] _122_\[21\] _06401_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__mux2_1
XFILLER_90_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12657_ _126_\[20\] _124_\[20\] _06368_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__mux2_1
XFILLER_128_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11608_ _05638_ _05640_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__nand2_1
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12588_ _06332_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11539_ _05558_ _05567_ _05568_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__a21o_1
XFILLER_116_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13209_ clknet_leaf_42_clk _00428_ VGND VGND VPWR VPWR _185_\[19\] sky130_fd_sc_hd__dfxtp_4
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08750_ _03136_ _03151_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__nor2_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08681_ _03105_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__xor2_4
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07701_ _02243_ _02244_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__nand2_1
XFILLER_93_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07632_ _01435_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__buf_2
XFILLER_81_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07563_ _01409_ _02111_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09302_ _03677_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__inv_2
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07494_ _02011_ _02038_ _02044_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__a21oi_1
X_06514_ _01214_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09233_ _02817_ _02787_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09164_ _185_\[23\] _03575_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__xnor2_1
X_08115_ _234_\[10\] _02564_ _02629_ _02635_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__a211o_1
XFILLER_135_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09095_ _170_\[21\] _02839_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__or2_1
X_08046_ _02577_ _02578_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__and2b_1
XFILLER_134_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09997_ _185_\[19\] _04150_ _04175_ _04375_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__o211a_1
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08948_ _03363_ _03365_ _03366_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__and3_1
XFILLER_91_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08879_ _03296_ _03299_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__xor2_1
XFILLER_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10910_ _04636_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__buf_2
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11890_ _140_\[0\] _140_\[2\] VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__xnor2_2
XFILLER_72_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10841_ _164_\[16\] _04983_ _05030_ _04998_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__o211a_1
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13560_ clknet_leaf_74_clk _00779_ VGND VGND VPWR VPWR _149_\[24\] sky130_fd_sc_hd__dfxtp_1
X_10772_ _173_\[29\] _04953_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__or2_1
X_13491_ clknet_leaf_46_clk _00710_ VGND VGND VPWR VPWR _158_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12511_ _06292_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12442_ _132_\[14\] _130_\[14\] _06247_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__mux2_1
XFILLER_40_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12373_ _06220_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11324_ _149_\[19\] _132_\[19\] VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__nand2_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11255_ _05327_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__and2_1
XFILLER_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10206_ _01239_ _04163_ _04416_ _04210_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__o31a_1
XFILLER_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11186_ _05267_ _05268_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__nor2_1
X_10137_ _04508_ _04509_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10068_ _04434_ _04443_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13827_ clknet_leaf_63_clk _01046_ VGND VGND VPWR VPWR _126_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13758_ clknet_leaf_57_clk _00977_ VGND VGND VPWR VPWR _132_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12709_ _124_\[13\] _122_\[13\] _06390_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__mux2_1
X_13689_ clknet_leaf_56_clk _00908_ VGND VGND VPWR VPWR _136_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09920_ _04011_ _04231_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__and2b_1
XFILLER_116_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09851_ _01283_ _03958_ _03904_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__o21a_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _142_\[9\] _04130_ _04131_ _04142_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_105_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08802_ _02037_ _03193_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__o21a_1
X_06994_ _243_\[28\] _01583_ _01557_ _01593_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__a211o_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08733_ _02846_ _03157_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__xnor2_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08664_ _02790_ _02845_ _02834_ _03091_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__o211a_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ _02160_ _02161_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08595_ _170_\[5\] _02784_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__or2_1
XFILLER_14_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07546_ _02066_ _02068_ _02093_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__and3_1
XFILLER_53_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07477_ _01428_ _02028_ _01495_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__a21oi_1
X_09216_ _03583_ _03585_ _03626_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__o21ba_1
XFILLER_108_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09147_ _228_\[22\] _231_\[22\] _03559_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__o21a_1
XFILLER_135_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09078_ _03491_ _03492_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__or2_1
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08029_ _02555_ _02556_ _02562_ _02355_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__a211o_1
XFILLER_123_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11040_ _04855_ _05164_ _05165_ _01436_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__a211o_1
XFILLER_131_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12991_ clknet_leaf_19_clk _00210_ VGND VGND VPWR VPWR _243_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11942_ _140_\[5\] _140_\[7\] VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11873_ _05864_ _05869_ _05867_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13612_ clknet_leaf_51_clk _00831_ VGND VGND VPWR VPWR _140_\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10824_ _170_\[12\] _05002_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__or2_1
X_13543_ clknet_leaf_73_clk _00762_ VGND VGND VPWR VPWR _149_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10755_ _173_\[24\] _04953_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__or2_1
X_10686_ _173_\[4\] _04917_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__or2_1
X_13474_ clknet_leaf_127_clk _00693_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfxtp_4
X_12425_ _06200_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__clkbuf_8
X_12356_ _06211_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11307_ _05279_ _05372_ _05373_ _05374_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__a31o_1
XFILLER_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12287_ _06174_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11238_ _05312_ _05313_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__nand2_1
XFILLER_106_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11169_ _05227_ _05254_ _05255_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__a21o_1
XFILLER_96_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07400_ _185_\[9\] _234_\[9\] VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__nand2_1
XFILLER_63_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08380_ _02827_ _02791_ _02824_ _02828_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__o211a_1
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07331_ _182_\[7\] _01626_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__nand2_1
XFILLER_35_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07262_ _01820_ _01821_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__nand2_1
XFILLER_117_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07193_ _01694_ _01754_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__xnor2_2
X_09001_ _03415_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__xor2_1
XFILLER_145_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09903_ _04277_ _04285_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__xor2_1
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09834_ _04209_ _04218_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__nor2_1
XFILLER_101_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _142_\[10\] _04152_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__and2_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06977_ _240_\[23\] _01565_ _01558_ _01581_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__o211a_1
X_09696_ _01241_ _01283_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__nor2_2
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08716_ _03101_ _03104_ _03141_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _185_\[6\] _03035_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__nand2_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _03004_ _03007_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__xnor2_4
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07529_ _02035_ _02052_ _02050_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__a21oi_1
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10540_ _173_\[21\] _04818_ _04820_ _04785_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__o211a_1
XFILLER_22_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10471_ _01225_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__buf_2
XFILLER_41_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12210_ _01393_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13190_ clknet_leaf_35_clk _00409_ VGND VGND VPWR VPWR _185_\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12141_ _140_\[31\] _142_\[31\] _06090_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__mux2_1
XFILLER_108_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12072_ _06049_ _06055_ _06060_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11023_ _03215_ _04630_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__nor2_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12974_ clknet_leaf_18_clk _00193_ VGND VGND VPWR VPWR _243_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11925_ _152_\[17\] _05914_ _05926_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__a21oi_1
XFILLER_72_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11856_ _05858_ _05860_ _05857_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__a21oi_2
XFILLER_33_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11787_ _05777_ _05783_ _05800_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__a21oi_1
X_10807_ _164_\[6\] _04986_ _05006_ _05001_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__a211o_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13526_ clknet_leaf_76_clk _00745_ VGND VGND VPWR VPWR _152_\[22\] sky130_fd_sc_hd__dfxtp_1
X_10738_ _167_\[18\] _04945_ _04957_ _04952_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__a211o_1
X_13457_ clknet_leaf_130_clk _00676_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_2
X_12408_ _06238_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__clkbuf_1
X_10669_ _176_\[31\] _04681_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__nor2_1
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13388_ clknet_leaf_12_clk _00607_ VGND VGND VPWR VPWR _167_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12339_ _06202_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06900_ _176_\[1\] _01523_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__or2_1
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07880_ _01684_ _01827_ _02178_ _02418_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__a211o_1
XFILLER_110_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06831_ _243_\[15\] _01474_ _01461_ _01475_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__o211a_1
XFILLER_95_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09550_ _03943_ _03944_ _03946_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__a21o_1
X_06762_ _01420_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__clkbuf_8
X_09481_ _195_\[3\] VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__clkinv_2
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08501_ _170_\[2\] _02776_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__nor2_1
X_06693_ _01378_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08432_ net59 _02868_ _01353_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__mux2_1
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08363_ _02002_ _02815_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__or2_1
X_07314_ _01840_ _01841_ _01871_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__a21o_1
X_08294_ _164_\[30\] _228_\[30\] _02750_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__mux2_1
X_07245_ _01654_ _01635_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07176_ _182_\[1\] _01604_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__nor2_1
XFILLER_133_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09817_ _04120_ _04145_ _04144_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__o21ai_1
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09748_ _04080_ _04107_ _04050_ _03872_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__o211a_1
XFILLER_100_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _03870_ _04070_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__nand2_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _118_\[5\] _118_\[16\] VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__xor2_1
XFILLER_70_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _124_\[4\] _122_\[4\] _06379_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__mux2_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _118_\[26\] _118_\[30\] VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__xnor2_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11572_ _118_\[23\] _118_\[2\] VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10523_ _173_\[16\] _04774_ _04808_ _04777_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__a211o_1
X_13311_ clknet_leaf_8_clk _00530_ VGND VGND VPWR VPWR _176_\[25\] sky130_fd_sc_hd__dfxtp_1
Xinput19 din[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10454_ _176_\[28\] _04725_ _04759_ _04728_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__a211o_1
X_13242_ clknet_leaf_6_clk _00461_ VGND VGND VPWR VPWR _182_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10385_ _179_\[9\] _182_\[9\] _04693_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__mux2_1
X_13173_ clknet_leaf_103_clk _00392_ VGND VGND VPWR VPWR _225_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12124_ _140_\[23\] _142_\[23\] _06079_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__mux2_1
XFILLER_78_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12055_ _142_\[29\] _06045_ _06005_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__mux2_1
XFILLER_89_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11006_ _164_\[3\] _04678_ _02946_ _04686_ _04648_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__o221a_1
XFILLER_46_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12957_ clknet_leaf_21_clk _00176_ VGND VGND VPWR VPWR _246_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12888_ _093_ _01296_ _04060_ _06487_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__a22o_1
X_11908_ _142_\[16\] _05911_ _05893_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__mux2_1
X_11839_ _05815_ _05825_ _05827_ _05848_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__o31a_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13509_ clknet_leaf_60_clk _00728_ VGND VGND VPWR VPWR _152_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07030_ _173_\[5\] _01620_ _01617_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__mux2_1
XFILLER_142_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08981_ _03359_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__inv_2
XFILLER_96_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07932_ _02465_ _02467_ _02468_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__or3_1
XFILLER_96_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07863_ _02398_ _02400_ _02401_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__and3_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09602_ _03989_ _03991_ _03995_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06814_ _246_\[10\] _01407_ _01460_ _01463_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__a211o_1
XFILLER_68_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09533_ _03879_ _03928_ _03929_ _195_\[4\] VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__a31o_1
XFILLER_56_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07794_ _02305_ _02324_ _02333_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__and3_1
XFILLER_37_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06745_ _01404_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__buf_4
X_09464_ _03866_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__inv_2
X_06676_ _01369_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08415_ net54 _02855_ _01353_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__mux2_1
X_09395_ _03800_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__inv_2
X_08346_ _02801_ _02791_ _02760_ _02802_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__o211a_1
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08277_ _164_\[25\] _228_\[25\] _02750_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__mux2_1
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07228_ _243_\[3\] _240_\[3\] _01612_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__mux2_2
XFILLER_20_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07159_ _01269_ _01711_ _01712_ _01722_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__a31o_1
XFILLER_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10170_ _04437_ _03893_ _04540_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__or3_1
XFILLER_120_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13860_ clknet_leaf_63_clk _01079_ VGND VGND VPWR VPWR _124_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13791_ clknet_leaf_65_clk _01010_ VGND VGND VPWR VPWR _130_\[31\] sky130_fd_sc_hd__dfxtp_1
X_12811_ _122_\[30\] _120_\[30\] _01367_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__mux2_1
XFILLER_28_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12742_ _06413_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__clkbuf_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _126_\[28\] _124_\[28\] _06368_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__mux2_1
XFILLER_63_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11624_ _116_\[21\] _05654_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__nand2_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11555_ _116_\[14\] _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__nand2_1
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11486_ _05518_ _05523_ _05517_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__a21bo_1
X_10506_ _173_\[11\] _04774_ _04796_ _04777_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__a211o_1
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13225_ clknet_leaf_24_clk _00444_ VGND VGND VPWR VPWR _182_\[3\] sky130_fd_sc_hd__dfxtp_1
X_10437_ _179_\[23\] _04721_ _04705_ _04747_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__o211a_1
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10368_ _176_\[3\] _04683_ _04698_ _01419_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__a211o_1
X_13156_ clknet_leaf_111_clk _00375_ VGND VGND VPWR VPWR _225_\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12107_ _06080_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10299_ _01217_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__clkbuf_4
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ clknet_leaf_104_clk _00306_ VGND VGND VPWR VPWR _234_\[31\] sky130_fd_sc_hd__dfxtp_1
X_12038_ _05991_ _06027_ _06029_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__o21ai_1
XFILLER_111_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06530_ _01238_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__clkbuf_4
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08200_ _164_\[3\] _228_\[3\] _02687_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__mux2_1
XFILLER_119_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09180_ _03589_ _03590_ _01354_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__o21a_1
X_08131_ _167_\[15\] _02616_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__or2_1
X_08062_ _01635_ _01620_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07013_ _01435_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__buf_2
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08964_ _02830_ _02790_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07915_ _185_\[26\] _234_\[26\] VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__or2_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08895_ _185_\[15\] _03314_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07846_ _185_\[24\] _234_\[24\] VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__nand2_1
XFILLER_83_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07777_ _02316_ _02318_ _01408_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__a21oi_1
X_09516_ _03913_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__buf_2
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06728_ _118_\[27\] _116_\[27\] _01394_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__mux2_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09447_ _02598_ _03850_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06659_ _01253_ _01324_ _01325_ _01356_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__nand4_1
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09378_ _03783_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__inv_2
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08329_ _228_\[6\] _02771_ _02765_ _02789_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__o211a_1
XFILLER_138_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11340_ _149_\[21\] _132_\[21\] VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__nand2_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11271_ _05341_ _05342_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__nand2_1
X_13010_ clknet_leaf_14_clk _00229_ VGND VGND VPWR VPWR _240_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10222_ _04572_ _04568_ _04590_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__nor3_1
XFILLER_106_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10153_ _04517_ _04523_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__and2_1
XFILLER_48_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10084_ _04075_ _03960_ _04278_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13912_ clknet_leaf_91_clk _01131_ VGND VGND VPWR VPWR _122_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13843_ clknet_leaf_94_clk _01062_ VGND VGND VPWR VPWR _126_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13774_ clknet_leaf_84_clk _00993_ VGND VGND VPWR VPWR _130_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10986_ net55 _05110_ _05132_ _05122_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__a211o_1
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12725_ _06404_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12656_ _01392_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__buf_4
XFILLER_31_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11607_ _05639_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__inv_2
X_12587_ _128_\[19\] _126_\[19\] _06324_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__mux2_1
XFILLER_128_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11538_ _05576_ _05577_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__nand2_1
X_11469_ _118_\[24\] _118_\[13\] VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13208_ clknet_leaf_41_clk _00427_ VGND VGND VPWR VPWR _185_\[18\] sky130_fd_sc_hd__dfxtp_4
XFILLER_124_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13139_ clknet_leaf_118_clk _00358_ VGND VGND VPWR VPWR _228_\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ _185_\[19\] _234_\[19\] VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__nand2_1
XFILLER_78_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08680_ _01927_ _03073_ _03106_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__o21a_1
XFILLER_38_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07631_ _01657_ _01973_ _01886_ _02177_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__o211a_1
XFILLER_38_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07562_ _02108_ _02110_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__xnor2_2
XFILLER_65_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06513_ _01224_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09301_ _185_\[26\] _03676_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__nand2_1
X_07493_ _02040_ _02043_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__xor2_1
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09232_ _02383_ _03641_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__nand2_1
XFILLER_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09163_ _02852_ _03574_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08114_ _231_\[10\] _02611_ _01695_ _02634_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__o211a_1
X_09094_ _170_\[21\] _02839_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__nand2_1
XFILLER_134_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08045_ _02540_ _02542_ _02541_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__a21bo_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09996_ _03945_ _04373_ _04374_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__or3_1
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08947_ _03095_ _03099_ _03238_ _03364_ _03360_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__a2111o_1
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08878_ _03251_ _03241_ _03297_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__a31o_1
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07829_ _02329_ _02331_ _02367_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__and3_1
XFILLER_17_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10840_ _05028_ _05029_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__or2_1
XFILLER_71_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10771_ _01225_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__clkbuf_4
X_13490_ clknet_leaf_42_clk _00709_ VGND VGND VPWR VPWR _158_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12510_ _130_\[14\] _128_\[14\] _06291_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__mux2_1
X_12441_ _06255_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12372_ _132_\[12\] _134_\[12\] _06219_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__mux2_1
XFILLER_125_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11323_ _149_\[19\] _132_\[19\] VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__nor2_1
Xclkbuf_4_0_0_clk clknet_3_0_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_141_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11254_ _149_\[10\] _132_\[10\] VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__nand2_1
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10205_ _04437_ _04158_ _04360_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__or3_1
XFILLER_69_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11185_ _149_\[1\] _132_\[1\] VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__nor2_1
XFILLER_69_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10136_ _04488_ _04491_ _04486_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__a21o_1
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10067_ _04210_ _04435_ _04439_ _04442_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__a31o_1
XFILLER_35_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13826_ clknet_leaf_63_clk _01045_ VGND VGND VPWR VPWR _126_\[2\] sky130_fd_sc_hd__dfxtp_1
X_13757_ clknet_leaf_57_clk _00976_ VGND VGND VPWR VPWR _132_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10969_ _164_\[22\] _05107_ _05094_ _05120_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__o211a_1
XFILLER_16_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12708_ _06395_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__clkbuf_1
X_13688_ clknet_leaf_56_clk _00907_ VGND VGND VPWR VPWR _136_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12639_ _06359_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09850_ _03905_ _03981_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__and2_1
XFILLER_124_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _04155_ _04168_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08801_ _185_\[11\] _03192_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__nand2_1
X_06993_ _240_\[28\] _01565_ _01558_ _01592_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__o211a_1
XFILLER_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _02807_ _02768_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08663_ _01856_ _03069_ _03090_ _02355_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__a211o_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07614_ _243_\[16\] _240_\[16\] _01657_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__mux2_4
XFILLER_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08594_ _03001_ _03022_ _01354_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__o21ai_1
XFILLER_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07545_ _02066_ _02068_ _02093_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__a21oi_1
XFILLER_41_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_127_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_127_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_22_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07476_ _02026_ _02027_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__xor2_4
X_09215_ _03581_ _03582_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__and2b_1
XFILLER_22_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09146_ _228_\[22\] _231_\[22\] _02842_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__a21o_1
XFILLER_135_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09077_ _03481_ _03482_ _03490_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__and3_1
XFILLER_123_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08028_ _01778_ _02561_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__nor2_1
XFILLER_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09979_ _04356_ _04357_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__or2_1
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12990_ clknet_leaf_22_clk _00209_ VGND VGND VPWR VPWR _243_\[30\] sky130_fd_sc_hd__dfxtp_1
X_11941_ _05941_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11872_ _05876_ _05878_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__nand2_1
XFILLER_72_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13611_ clknet_leaf_52_clk _00830_ VGND VGND VPWR VPWR _140_\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_72_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_118_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_118_clk sky130_fd_sc_hd__clkbuf_16
X_10823_ _164_\[11\] _04983_ _05017_ _04998_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__o211a_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13542_ clknet_leaf_65_clk _00761_ VGND VGND VPWR VPWR _149_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10754_ _167_\[23\] _04925_ _04968_ _04939_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__o211a_1
XFILLER_9_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13473_ clknet_leaf_122_clk _00692_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfxtp_1
XFILLER_13_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10685_ _167_\[3\] _04836_ _04919_ _04914_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__a211o_1
XFILLER_145_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12424_ _06246_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__clkbuf_1
X_12355_ _132_\[4\] _134_\[4\] _06208_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__mux2_1
XFILLER_65_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11306_ _152_\[16\] _01368_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__and2_1
XFILLER_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12286_ _136_\[4\] _134_\[4\] _06167_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__mux2_1
XFILLER_114_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11237_ _149_\[8\] _132_\[8\] VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__nand2_1
X_11168_ net21 _05202_ _05192_ _158_\[19\] VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__a22o_1
XFILLER_110_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10119_ _185_\[24\] _03867_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__or2_1
X_11099_ _158_\[1\] _158_\[0\] _158_\[2\] VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__nor3_1
XFILLER_82_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_109_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_109_clk sky130_fd_sc_hd__clkbuf_16
X_13809_ clknet_leaf_95_clk _01028_ VGND VGND VPWR VPWR _128_\[17\] sky130_fd_sc_hd__dfxtp_1
X_07330_ _182_\[7\] _01626_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__or2_1
XFILLER_16_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07261_ _182_\[4\] _01616_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__nand2_1
X_09000_ _02205_ _03384_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__o21a_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_07192_ _01645_ _01629_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09902_ _01232_ _04279_ _04281_ _04282_ _04284_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__a32o_1
XFILLER_116_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09833_ _04209_ _04218_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__and2_1
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09764_ _246_\[10\] _01314_ _03914_ _243_\[10\] _01462_ VGND VGND VPWR VPWR _04152_
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06976_ _176_\[23\] _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__or2_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09695_ _01235_ _03875_ _04005_ _04085_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__or4_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08715_ _185_\[8\] _03103_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__nand2_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _01927_ _03073_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__xnor2_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _185_\[5\] _03006_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__xnor2_4
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07528_ _02076_ _02077_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__and2b_1
X_07459_ _185_\[11\] _234_\[11\] VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__nand2_1
X_10470_ _173_\[1\] _04735_ _04770_ _04740_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__o211a_1
XFILLER_10_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09129_ _03468_ _03508_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__nand2_1
XFILLER_136_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12140_ _06097_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12071_ _140_\[18\] _06059_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11022_ net37 _04848_ _05153_ _05122_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__a211o_1
XFILLER_131_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12973_ clknet_leaf_19_clk _00192_ VGND VGND VPWR VPWR _243_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11924_ _152_\[17\] _05914_ _05903_ _152_\[16\] VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__o211a_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11855_ _05863_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__clkbuf_1
X_11786_ _05780_ _05792_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__nand2_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10806_ _167_\[6\] _04980_ _04958_ _05005_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__o211a_1
XFILLER_13_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13525_ clknet_leaf_78_clk _00744_ VGND VGND VPWR VPWR _152_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10737_ _170_\[18\] _04942_ _04922_ _04956_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__o211a_1
X_13456_ clknet_leaf_1_clk _00675_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_4
X_12407_ _132_\[29\] _134_\[29\] _06230_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__mux2_1
X_10668_ _173_\[31\] _04848_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__nand2_1
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13387_ clknet_leaf_12_clk _00606_ VGND VGND VPWR VPWR _167_\[5\] sky130_fd_sc_hd__dfxtp_1
X_10599_ _04724_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__buf_6
X_12338_ _136_\[28\] _134_\[28\] _06201_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__mux2_1
XFILLER_5_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12269_ _138_\[28\] _136_\[28\] _06156_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__mux2_1
XFILLER_99_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06830_ _179_\[15\] _01300_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__or2_1
XFILLER_95_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06761_ _01411_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__clkbuf_4
X_09480_ _03877_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__buf_4
X_06692_ _118_\[11\] _116_\[11\] _01370_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__mux2_1
X_08500_ _170_\[2\] _02776_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__and2_1
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08431_ _225_\[30\] VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__buf_4
XFILLER_36_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08362_ net41 _02814_ _01353_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__mux2_1
X_07313_ _01867_ _01870_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__xor2_1
X_08293_ _231_\[29\] _02730_ _02753_ _02762_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__a211o_1
X_07244_ _01781_ _01782_ _01783_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__nand3_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07175_ _182_\[1\] _01604_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__and2_1
XFILLER_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09816_ _04122_ _04147_ _04201_ _04124_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__or4b_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09747_ _04056_ _04135_ _01231_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__a21oi_1
X_06959_ _01518_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__buf_4
XFILLER_74_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09678_ _04066_ _04069_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__xnor2_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _02940_ _02974_ _02975_ _03057_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__a31o_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11640_ _05669_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__clkbuf_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11571_ _05607_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10522_ _176_\[16\] _04771_ _04806_ _04807_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__o211a_1
X_13310_ clknet_leaf_8_clk _00529_ VGND VGND VPWR VPWR _176_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13241_ clknet_leaf_6_clk _00460_ VGND VGND VPWR VPWR _182_\[19\] sky130_fd_sc_hd__dfxtp_1
X_10453_ _179_\[28\] _04721_ _04751_ _04758_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__o211a_1
XFILLER_6_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10384_ _176_\[8\] _04683_ _04709_ _01419_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__a211o_1
X_13172_ clknet_leaf_104_clk _00391_ VGND VGND VPWR VPWR _225_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12123_ _06088_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12054_ net22 _06044_ _05785_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__mux2_1
XFILLER_96_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11005_ net58 _04849_ _05144_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__a21o_1
XFILLER_93_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12956_ clknet_leaf_21_clk _00175_ VGND VGND VPWR VPWR _246_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12887_ _06489_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__clkbuf_1
X_11907_ net8 _05910_ _05852_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__mux2_1
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11838_ _05823_ _05835_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__and2_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13508_ clknet_leaf_58_clk _00727_ VGND VGND VPWR VPWR _152_\[4\] sky130_fd_sc_hd__dfxtp_1
X_11769_ _01358_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_40_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_127_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13439_ clknet_leaf_126_clk _00658_ VGND VGND VPWR VPWR _164_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08980_ _03395_ _03397_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__nand2_1
XFILLER_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07931_ _02394_ _02433_ _02435_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07862_ _02144_ _02147_ _02277_ _02399_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__a211o_1
X_09601_ _03988_ _03973_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__and2b_1
X_06813_ _243_\[10\] _01438_ _01461_ _01462_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__o211a_1
XFILLER_96_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09532_ _03874_ _195_\[0\] _01279_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__or3b_2
XFILLER_113_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07793_ _02305_ _02324_ _02333_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__a21oi_1
X_06744_ _01321_ _01358_ _01403_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__nor3_4
XFILLER_64_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06675_ _118_\[3\] _116_\[3\] _01368_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__mux2_1
X_09463_ _01418_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__buf_6
X_09394_ _03756_ _03777_ _03799_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__o21ai_1
X_08414_ _225_\[26\] VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__buf_6
XFILLER_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08345_ net37 _02798_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_31_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_137_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08276_ _01518_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__buf_4
X_07227_ _01786_ _01787_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__or2_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07158_ _01720_ _01721_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__nor2_1
XFILLER_133_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07089_ _240_\[18\] _01649_ _01607_ _01666_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__a211o_1
XFILLER_78_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_98_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_59_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12810_ _06448_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13790_ clknet_leaf_65_clk _01009_ VGND VGND VPWR VPWR _130_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12741_ _124_\[28\] _122_\[28\] _06412_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__mux2_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12672_ _06376_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11623_ _118_\[7\] _05653_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__xnor2_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11554_ _118_\[21\] _05591_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11485_ _05528_ _05529_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__or2b_1
X_10505_ _176_\[11\] _04771_ _04751_ _04795_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__o211a_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13224_ clknet_leaf_28_clk _00443_ VGND VGND VPWR VPWR _182_\[2\] sky130_fd_sc_hd__dfxtp_1
X_10436_ _182_\[23\] _04746_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__or2_1
XFILLER_124_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10367_ _179_\[3\] _04684_ _04686_ _04697_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__o211a_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13155_ clknet_leaf_112_clk _00374_ VGND VGND VPWR VPWR _225_\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12106_ _140_\[14\] _142_\[14\] _06079_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__mux2_1
XFILLER_105_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10298_ _179_\[10\] _04629_ _04653_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__a21o_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13086_ clknet_leaf_104_clk _00305_ VGND VGND VPWR VPWR _234_\[30\] sky130_fd_sc_hd__dfxtp_1
X_12037_ _06010_ _06013_ _06022_ _06028_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_89_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_78_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12939_ clknet_leaf_21_clk _00158_ VGND VGND VPWR VPWR _246_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08130_ _01406_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08061_ _02580_ _02582_ _02579_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07012_ _240_\[1\] _01601_ _01598_ _01606_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__o211a_1
XFILLER_143_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08963_ _03354_ _03356_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__and2b_1
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07914_ _01667_ _02450_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__xnor2_4
XFILLER_111_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08894_ _02862_ _03313_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07845_ _185_\[24\] _234_\[24\] VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__or2_1
XFILLER_140_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07776_ _02275_ _02281_ _02317_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__a21bo_1
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09515_ _392_\[4\] _01206_ _01246_ _01268_ _01251_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__o32ai_4
X_06727_ _01397_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__clkbuf_1
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09446_ _03847_ _03849_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06658_ _099_ _01328_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__nand2_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06589_ _01284_ _01276_ _01281_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__a21oi_1
XFILLER_12_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09377_ _03781_ _03782_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__nand2_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08328_ _02749_ _02788_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__or2_1
X_08259_ _231_\[19\] _02730_ _02712_ _02738_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__a211o_1
XFILLER_119_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11270_ _149_\[12\] _132_\[12\] VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__nand2_1
X_10221_ _04588_ _04589_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__or2b_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10152_ _04517_ _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__nor2_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10083_ _01281_ _03934_ _03904_ _03905_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__o22a_1
XFILLER_102_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13911_ clknet_leaf_92_clk _01130_ VGND VGND VPWR VPWR _122_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13842_ clknet_leaf_94_clk _01061_ VGND VGND VPWR VPWR _126_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13773_ clknet_leaf_84_clk _00992_ VGND VGND VPWR VPWR _130_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10985_ _164_\[27\] _05107_ _04865_ _05131_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__o211a_1
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12724_ _124_\[20\] _122_\[20\] _06401_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__mux2_1
XFILLER_43_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12655_ _06367_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11606_ _116_\[19\] _05637_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__nor2_1
X_12586_ _06331_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11537_ _116_\[12\] _05575_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__or2_1
XFILLER_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11468_ _05514_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11399_ _05453_ _05454_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__nand2_1
X_13207_ clknet_leaf_42_clk _00426_ VGND VGND VPWR VPWR _185_\[17\] sky130_fd_sc_hd__dfxtp_4
X_10419_ _176_\[18\] _04691_ _04734_ _04677_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__o211a_1
XFILLER_124_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13138_ clknet_leaf_118_clk _00357_ VGND VGND VPWR VPWR _228_\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ clknet_leaf_83_clk _00288_ VGND VGND VPWR VPWR _234_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_66_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07630_ _01355_ _02166_ _02167_ _02176_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__a31o_1
XFILLER_54_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07561_ _02056_ _02109_ _02081_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__o21ai_2
XFILLER_65_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06512_ _01222_ _01223_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__and2_1
X_09300_ _02460_ _03681_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__nand2_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07492_ _02041_ _02042_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__nand2_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09231_ _03613_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__inv_2
X_09162_ _02811_ _02781_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08113_ _167_\[10\] _02616_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__or2_1
X_09093_ _02835_ _01426_ _03379_ _03507_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__o211a_1
X_08044_ _02573_ _02576_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09995_ _04345_ _04352_ _04372_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__a21oi_1
XFILLER_103_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08946_ _03239_ _03364_ _03360_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__or3_1
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08877_ _03252_ _03266_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__nor2_1
XFILLER_28_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07828_ _02329_ _02331_ _02367_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__a21oi_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07759_ _02270_ _02271_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__and2b_1
XFILLER_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10770_ _167_\[28\] _04925_ _04979_ _04939_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__o211a_1
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09429_ _03832_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__nand2_1
X_12440_ _132_\[13\] _130_\[13\] _06247_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__mux2_1
XFILLER_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12371_ _06004_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__clkbuf_4
XFILLER_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11322_ _05279_ _05385_ _05386_ _05387_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__a31o_1
XFILLER_134_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11253_ _149_\[10\] _132_\[10\] VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__or2_1
X_10204_ _04560_ _04564_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__nor2_1
XFILLER_106_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11184_ _149_\[1\] _132_\[1\] VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__and2_1
XFILLER_122_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10135_ _04505_ _04507_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__nand2_1
XFILLER_67_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10066_ _01238_ _04440_ _04441_ _01232_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__o211a_1
XFILLER_85_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13825_ clknet_leaf_64_clk _01044_ VGND VGND VPWR VPWR _126_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13756_ clknet_leaf_67_clk _00975_ VGND VGND VPWR VPWR _132_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10968_ _167_\[22\] _05089_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__or2_1
X_13687_ clknet_leaf_67_clk _00906_ VGND VGND VPWR VPWR _136_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12707_ _124_\[12\] _122_\[12\] _06390_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__mux2_1
X_10899_ _05028_ _05071_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__or2_1
X_12638_ _126_\[11\] _124_\[11\] _06357_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__mux2_1
XFILLER_129_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12569_ _06322_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08800_ _02071_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__xnor2_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09780_ _04159_ _04162_ _04167_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__and3_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06992_ _176_\[28\] _01580_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__or2_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _02797_ _03032_ _02861_ _03156_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__a211o_1
X_08662_ _01923_ _03089_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__nor2_1
XFILLER_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07613_ _02158_ _02159_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__or2_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08593_ _03001_ _03022_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__and2_1
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07544_ _02089_ _02092_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__xor2_1
X_07475_ _01998_ _02000_ _01996_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__o21a_2
XFILLER_50_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09214_ _03622_ _03624_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__xnor2_1
X_09145_ _03555_ _03557_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__xor2_1
XFILLER_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09076_ _03481_ _03482_ _03490_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__a21oi_1
X_08027_ _02559_ _02560_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__xnor2_2
XFILLER_116_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09978_ _04354_ _04355_ _142_\[19\] VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__a21oi_1
XFILLER_76_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08929_ _03341_ _03342_ _03346_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__nand3_1
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11940_ _142_\[19\] _05940_ _05893_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__mux2_1
XFILLER_85_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11871_ _05877_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__inv_2
XFILLER_84_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13610_ clknet_leaf_52_clk _00829_ VGND VGND VPWR VPWR _140_\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10822_ _04971_ _05016_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__or2_1
X_13541_ clknet_leaf_63_clk _00760_ VGND VGND VPWR VPWR _149_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10753_ _04888_ _04967_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__or2_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10684_ _170_\[3\] _04833_ _04806_ _04918_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__o211a_1
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13472_ clknet_leaf_122_clk _00691_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfxtp_4
XFILLER_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12423_ _132_\[5\] _130_\[5\] _06201_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__mux2_1
X_12354_ _06210_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11305_ _05355_ _05364_ _05361_ _05370_ _05360_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__a311o_1
XFILLER_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12285_ _06173_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11236_ _149_\[8\] _132_\[8\] VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__or2_1
XFILLER_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11167_ _158_\[19\] _01264_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10118_ _04488_ _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__xor2_1
XFILLER_110_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11098_ _05190_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__buf_2
X_10049_ _04379_ _04390_ _04424_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__or3_1
XFILLER_48_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13808_ clknet_leaf_95_clk _01027_ VGND VGND VPWR VPWR _128_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13739_ clknet_leaf_48_clk _00958_ VGND VGND VPWR VPWR _132_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07260_ _182_\[4\] _01616_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__or2_1
X_07191_ _01733_ _01734_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__and2b_1
XFILLER_145_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09901_ _01231_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__nor2_1
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09832_ _04210_ _04212_ _04213_ _04217_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__a31o_1
XFILLER_101_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09763_ _04128_ _04146_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__nand2_1
XFILLER_112_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08714_ _01974_ _03139_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__xnor2_1
X_06975_ _01339_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__clkbuf_2
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _03884_ _03927_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__nand2_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08645_ _185_\[7\] _03072_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08576_ _02858_ _03005_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__xnor2_4
X_07527_ _02045_ _02061_ _02075_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__or3_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07458_ _185_\[11\] _234_\[11\] VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__or2_1
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07389_ _01923_ _01944_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__nor2_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09128_ _03539_ _03540_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__nor2_1
XFILLER_135_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09059_ _170_\[19\] _02830_ _03472_ _03473_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__a211oi_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12070_ _140_\[16\] _152_\[31\] VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11021_ _03184_ _04865_ _164_\[10\] _04684_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_131_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12972_ clknet_leaf_17_clk _00191_ VGND VGND VPWR VPWR _243_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11923_ _05906_ _05915_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__or2_1
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11854_ _142_\[11\] _05862_ _05765_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__mux2_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10805_ _170_\[6\] _05002_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__or2_1
X_11785_ _05799_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13524_ clknet_leaf_75_clk _00743_ VGND VGND VPWR VPWR _152_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10736_ _173_\[18\] _04953_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__or2_1
X_10667_ _02570_ _04861_ _04906_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__a21o_1
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13455_ clknet_leaf_113_clk _00674_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_4
X_12406_ _06237_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10598_ _173_\[7\] _04629_ _04860_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__o21a_1
X_13386_ clknet_leaf_11_clk _00605_ VGND VGND VPWR VPWR _167_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12337_ _06200_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__clkbuf_4
X_12268_ _06164_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__clkbuf_1
X_11219_ _152_\[5\] _05297_ _01362_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__mux2_1
X_12199_ _06128_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06760_ _246_\[0\] _01407_ _01414_ _01419_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__a211o_1
XFILLER_55_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06691_ _01377_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08430_ _228_\[29\] _02838_ _02861_ _02867_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__a211o_1
XFILLER_36_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08361_ _225_\[14\] VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__clkbuf_4
X_07312_ _01868_ _01869_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__nand2_1
X_08292_ _228_\[29\] _02733_ _02760_ _02761_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__o211a_1
X_07243_ _01788_ _01789_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__and2b_1
XFILLER_20_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07174_ _01720_ _01735_ _01518_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09815_ _04171_ _04194_ _04195_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__nand3_1
XFILLER_113_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09746_ _01242_ _03890_ _03898_ _03872_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__a31oi_1
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06958_ _01405_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__clkbuf_2
XFILLER_74_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09677_ _04067_ _04068_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__or2_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06889_ _01302_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__buf_4
X_08628_ _02973_ _03026_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__nand2_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _02987_ _02989_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11570_ _149_\[15\] _05606_ _05533_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__mux2_1
XFILLER_23_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10521_ _179_\[16\] _04799_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__or2_1
XFILLER_50_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13240_ clknet_leaf_25_clk _00459_ VGND VGND VPWR VPWR _182_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10452_ _182_\[28\] _04746_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__or2_1
X_10383_ _179_\[8\] _04684_ _04705_ _04708_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__o211a_1
X_13171_ clknet_leaf_105_clk _00390_ VGND VGND VPWR VPWR _225_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12122_ _140_\[22\] _142_\[22\] _06079_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__mux2_1
XFILLER_123_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12053_ _06038_ _06043_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11004_ _164_\[2\] net68 _02936_ _04692_ _01417_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__a221o_1
XFILLER_131_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_77_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12955_ clknet_leaf_21_clk _00174_ VGND VGND VPWR VPWR _246_\[27\] sky130_fd_sc_hd__dfxtp_1
X_11906_ _05906_ _05909_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__xor2_1
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12886_ _03864_ _06488_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__and2_1
XFILLER_73_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11837_ _05845_ _05846_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__nand2_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11768_ _05777_ _05783_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__or2_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ clknet_leaf_60_clk _00726_ VGND VGND VPWR VPWR _152_\[3\] sky130_fd_sc_hd__dfxtp_1
X_10719_ _170_\[13\] _04942_ _04922_ _04943_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__o211a_1
X_11699_ _118_\[4\] _118_\[15\] VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__or2_1
XFILLER_127_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13438_ clknet_leaf_126_clk _00657_ VGND VGND VPWR VPWR _164_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13369_ clknet_leaf_125_clk _00588_ VGND VGND VPWR VPWR _170_\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07930_ _02402_ _02466_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__nor2_1
XFILLER_122_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07861_ _02280_ _02399_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__or2_1
X_09600_ _185_\[3\] _03869_ _03919_ _03994_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__o211a_1
XFILLER_110_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06812_ _179_\[10\] _01300_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__or2_1
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07792_ _02331_ _02332_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__nand2_1
X_09531_ _01279_ _195_\[0\] _03874_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__or3b_4
X_06743_ _01323_ _01307_ _01304_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__a21oi_2
XFILLER_110_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06674_ _01367_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__buf_4
XFILLER_64_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09462_ _03859_ _03863_ _03865_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09393_ _03796_ _03798_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__xnor2_1
X_08413_ _228_\[25\] _02838_ _02810_ _02854_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__a211o_1
X_08344_ _225_\[10\] VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08275_ _01404_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__buf_2
XFILLER_20_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07226_ _01756_ _01779_ _01785_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__and3_1
X_07157_ _01718_ _01719_ _01302_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__o21ai_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07088_ _01664_ _01639_ _01609_ _01665_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__o211a_1
XFILLER_120_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09729_ _04117_ _04118_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__nor2_1
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12740_ _01392_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__clkbuf_4
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12671_ _126_\[27\] _124_\[27\] _06368_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__mux2_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11622_ _118_\[24\] _118_\[28\] VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__xnor2_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11553_ _118_\[17\] _118_\[0\] VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11484_ _116_\[7\] _05527_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__nand2_1
X_10504_ _179_\[11\] _04746_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__or2_1
X_13223_ clknet_leaf_28_clk _00442_ VGND VGND VPWR VPWR _182_\[1\] sky130_fd_sc_hd__dfxtp_2
X_10435_ _01216_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__buf_2
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13154_ clknet_leaf_2_clk _00373_ VGND VGND VPWR VPWR _225_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12105_ _06004_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__clkbuf_4
X_10366_ _182_\[3\] _04696_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__or2_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10297_ _182_\[10\] _01218_ _04642_ _04650_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__a31o_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13085_ clknet_leaf_102_clk _00304_ VGND VGND VPWR VPWR _234_\[29\] sky130_fd_sc_hd__dfxtp_1
X_12036_ _06008_ _06021_ _06020_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__o21ba_1
XFILLER_111_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12938_ clknet_leaf_21_clk _00157_ VGND VGND VPWR VPWR _246_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _06479_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ _02585_ _02588_ _02584_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__o21bai_1
XFILLER_127_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07011_ _01568_ _01605_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__or2_1
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08962_ _03351_ _03353_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__nor2_1
XFILLER_130_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07913_ _01620_ _237_\[0\] VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__xnor2_2
XFILLER_69_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08893_ _02823_ _02784_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07844_ _01704_ _02382_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__xnor2_4
XFILLER_57_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07775_ _02274_ _02272_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__or2b_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09514_ _03871_ _03882_ _03895_ _03911_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__a31o_1
X_06726_ _118_\[26\] _116_\[26\] _01394_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__mux2_1
X_06657_ _01266_ _01355_ _01211_ VGND VGND VPWR VPWR _436_\[4\] sky130_fd_sc_hd__o21ai_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09445_ _02871_ _231_\[31\] _03848_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__o21a_1
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06588_ _01276_ _01285_ _01293_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__a21oi_1
XFILLER_40_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09376_ _185_\[29\] _03780_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__or2_1
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08327_ net64 _02787_ _02750_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__mux2_1
X_08258_ _228_\[19\] _02733_ _02723_ _02737_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__o211a_1
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07209_ _01710_ _01770_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__or2_1
X_10220_ _04558_ _04573_ _04587_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__or3b_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08189_ _164_\[0\] _228_\[0\] _02687_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__mux2_1
X_10151_ _01239_ _04519_ _04522_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__a21o_1
XFILLER_106_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10082_ _04060_ _03984_ _04025_ _04418_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__and4_1
XFILLER_121_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13910_ clknet_leaf_96_clk _01129_ VGND VGND VPWR VPWR _122_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13841_ clknet_leaf_95_clk _01060_ VGND VGND VPWR VPWR _126_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13772_ clknet_leaf_87_clk _00991_ VGND VGND VPWR VPWR _130_\[12\] sky130_fd_sc_hd__dfxtp_1
X_10984_ _167_\[27\] _04867_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__or2_1
XFILLER_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12723_ _06403_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12654_ _126_\[19\] _124_\[19\] _06357_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__mux2_1
XFILLER_30_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11605_ _116_\[19\] _05637_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__nand2_1
X_12585_ _128_\[18\] _126_\[18\] _06324_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__mux2_1
XFILLER_129_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11536_ _116_\[12\] _05575_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__nand2_1
XFILLER_137_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11467_ _149_\[5\] _05513_ _05439_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__mux2_1
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13206_ clknet_leaf_41_clk _00425_ VGND VGND VPWR VPWR _185_\[16\] sky130_fd_sc_hd__dfxtp_2
X_11398_ _149_\[28\] _132_\[28\] VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__or2_1
X_10418_ _04712_ _04733_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__or2_1
XFILLER_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10349_ _04682_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__buf_4
XFILLER_3_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13137_ clknet_leaf_118_clk _00356_ VGND VGND VPWR VPWR _228_\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13068_ clknet_leaf_83_clk _00287_ VGND VGND VPWR VPWR _234_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _05984_ _05998_ _06012_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__o21a_1
XFILLER_120_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07560_ _182_\[13\] _01645_ _01642_ _182_\[12\] VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__a22o_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06511_ _190_\[1\] _190_\[0\] _01215_ _190_\[2\] VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__a31o_1
XFILLER_62_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07491_ _185_\[12\] _234_\[12\] VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__nand2_1
X_09230_ _185_\[24\] _03612_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__nand2_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09161_ _185_\[22\] _03548_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__nand2_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08112_ _234_\[9\] _02448_ _02419_ _02633_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__o211a_1
X_09092_ _01856_ _03478_ _03506_ _01495_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__a211o_1
XFILLER_30_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08043_ _02574_ _02575_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__nor2_1
XFILLER_134_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09994_ _04345_ _04352_ _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__and3_1
XFILLER_103_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08945_ _03236_ _03267_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__nand2_1
XFILLER_111_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08876_ _03252_ _03266_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__nand2_1
XFILLER_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07827_ _02365_ _02366_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__nand2_1
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07758_ _02298_ _02299_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__xnor2_4
X_06709_ _118_\[19\] _116_\[19\] _01381_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__mux2_1
XFILLER_25_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07689_ _182_\[19\] _01667_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__nor2_1
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09428_ _03794_ _03813_ _03831_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__or3_1
XFILLER_9_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09359_ _03764_ _03739_ _03740_ _01923_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__a31oi_1
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12370_ _06218_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11321_ _152_\[18\] _01368_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__and2_1
XFILLER_125_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11252_ _05326_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11183_ _152_\[0\] _05262_ _05266_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__a21o_1
X_10203_ _04565_ _04566_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__nor2_1
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10134_ _04506_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__inv_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10065_ _03873_ _03876_ _04027_ _04303_ _04078_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__a2111o_1
XFILLER_125_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13824_ clknet_leaf_64_clk _01043_ VGND VGND VPWR VPWR _126_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13755_ clknet_leaf_57_clk _00974_ VGND VGND VPWR VPWR _132_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10967_ net49 _05110_ _05119_ _05086_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__a211o_1
X_13686_ clknet_leaf_56_clk _00905_ VGND VGND VPWR VPWR _136_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10898_ _164_\[1\] _167_\[1\] _05064_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__mux2_1
X_12706_ _06394_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__clkbuf_1
X_12637_ _06358_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12568_ _128_\[10\] _126_\[10\] _06313_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__mux2_1
X_12499_ _130_\[9\] _128_\[9\] _06280_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__mux2_1
XFILLER_129_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11519_ _05542_ _05549_ _05550_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__a21o_1
XFILLER_109_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06991_ _243_\[27\] _01583_ _01557_ _01591_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__a211o_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _01520_ _03133_ _03155_ _02202_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__o211a_1
XFILLER_94_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08661_ _03086_ _03088_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07612_ _02119_ _02121_ _02157_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__and3_1
XFILLER_54_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08592_ _03020_ _03021_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__or2b_1
XFILLER_81_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07543_ _02090_ _02091_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__nand2_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07474_ _02024_ _02025_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__nand2_2
XFILLER_50_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09213_ _228_\[24\] _231_\[24\] _03623_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__o21a_1
XFILLER_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09144_ _02311_ _03526_ _03556_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__a21o_1
XFILLER_108_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09075_ _02271_ _03489_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08026_ _02531_ _02532_ _02533_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__o21a_1
XFILLER_89_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09977_ _142_\[19\] _04354_ _04355_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__and3_1
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08928_ _03341_ _03342_ _03346_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__a21o_1
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08859_ _185_\[14\] _03279_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11870_ _152_\[13\] _05875_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__nor2_1
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10821_ _167_\[11\] _170_\[11\] _04995_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__mux2_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13540_ clknet_leaf_65_clk _00759_ VGND VGND VPWR VPWR _149_\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10752_ _170_\[23\] _173_\[23\] _04936_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__mux2_1
XFILLER_13_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13471_ clknet_leaf_122_clk _00690_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfxtp_4
XFILLER_13_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12422_ _06245_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__clkbuf_1
X_10683_ _173_\[3\] _04917_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__or2_1
XFILLER_9_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12353_ _132_\[3\] _134_\[3\] _06208_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__mux2_1
XFILLER_138_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12284_ _136_\[3\] _134_\[3\] _06167_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__mux2_1
X_11304_ _05370_ _05371_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__nand2_1
X_11235_ _05311_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11166_ _05227_ _05252_ _05253_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__a21o_1
X_11097_ _05199_ _05197_ _05200_ _05201_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__o22ai_1
X_10117_ _04451_ _04452_ _04489_ _04490_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__o31a_1
XFILLER_110_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10048_ _04379_ _04390_ _04424_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__o21a_1
XFILLER_48_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13807_ clknet_leaf_98_clk _01026_ VGND VGND VPWR VPWR _128_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11999_ _05994_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__clkbuf_1
X_13738_ clknet_leaf_77_clk _00957_ VGND VGND VPWR VPWR _132_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13669_ clknet_leaf_59_clk _00888_ VGND VGND VPWR VPWR _136_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07190_ _01731_ _01732_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__nor2_1
XFILLER_144_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09900_ _03886_ _03907_ _04139_ _01237_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__o211a_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09831_ _01236_ _04214_ _04216_ _03871_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__o211a_1
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _03868_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__buf_2
XFILLER_112_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06974_ _243_\[22\] _01548_ _01545_ _01579_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__o211a_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08713_ _185_\[9\] _03138_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__xnor2_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _04075_ _04080_ _04083_ _03872_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__a211o_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08644_ _02865_ _03071_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__xnor2_2
XFILLER_82_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08575_ _02827_ _02790_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__xnor2_2
XFILLER_81_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07526_ _02045_ _02061_ _02075_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__o21a_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07457_ _01678_ _02008_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07388_ _01924_ _01925_ _01943_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__o21a_1
XFILLER_10_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09127_ _170_\[22\] _02842_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__and2_1
XFILLER_135_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09058_ _170_\[19\] _02830_ _03435_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__o21a_1
XFILLER_135_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08009_ _02541_ _02542_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__nand2_1
XFILLER_135_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11020_ net67 _04849_ _05152_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__a21o_1
XFILLER_77_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12971_ clknet_leaf_18_clk _00190_ VGND VGND VPWR VPWR _243_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11922_ _05922_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__nand2_1
X_11853_ net3 _05861_ _05852_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__mux2_1
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10804_ _164_\[5\] _04986_ _05004_ _05001_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__a211o_1
XFILLER_14_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11784_ _142_\[5\] _05798_ _05765_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__mux2_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13523_ clknet_leaf_78_clk _00742_ VGND VGND VPWR VPWR _152_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10735_ _167_\[17\] _04945_ _04955_ _04952_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__a211o_1
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10666_ _176_\[30\] net68 _04638_ _173_\[30\] _02711_ VGND VGND VPWR VPWR _04906_
+ sky130_fd_sc_hd__a221o_1
X_13454_ clknet_leaf_113_clk _00673_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfxtp_4
XFILLER_127_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12405_ _132_\[28\] _134_\[28\] _06230_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__mux2_1
XFILLER_9_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13385_ clknet_leaf_1_clk _00604_ VGND VGND VPWR VPWR _167_\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10597_ _176_\[7\] _04678_ _01892_ _04686_ _04648_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__o221a_1
XFILLER_114_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12336_ _01366_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__buf_4
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12267_ _138_\[27\] _136_\[27\] _06156_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__mux2_1
X_11218_ _05295_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__xnor2_1
X_12198_ _140_\[26\] _138_\[26\] _06123_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__mux2_1
XFILLER_96_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11149_ net16 _05202_ _05193_ _158_\[14\] VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__a22o_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06690_ _118_\[10\] _116_\[10\] _01370_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__mux2_1
X_08360_ _228_\[13\] _02775_ _02810_ _02813_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__a211o_1
X_07311_ _185_\[6\] _234_\[6\] VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__or2_1
XFILLER_32_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08291_ _164_\[29\] _02736_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__or2_1
XFILLER_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07242_ _01794_ _01796_ _01793_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07173_ _01720_ _01735_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__and2_1
XFILLER_145_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09814_ _185_\[11\] _04150_ _04175_ _04200_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__o211a_1
XFILLER_98_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09745_ _03886_ _04010_ _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__or3_1
X_06957_ _243_\[17\] _01536_ _01557_ _01567_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__a211o_1
X_09676_ _03996_ _04018_ _04039_ _04040_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__o211a_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ _246_\[30\] _01496_ _01509_ _01517_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__a211o_1
XFILLER_39_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08627_ _03054_ _03055_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__nand2_1
XFILLER_27_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _01789_ _02956_ _02988_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__a21oi_1
X_07509_ _01884_ _02059_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__nor2_1
X_08489_ _02919_ _02921_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10520_ _04685_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__buf_2
XFILLER_109_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10451_ _176_\[27\] _04725_ _04757_ _04728_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__a211o_1
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10382_ _182_\[8\] _04696_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__or2_1
X_13170_ clknet_leaf_100_clk _00389_ VGND VGND VPWR VPWR _225_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12121_ _06087_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12052_ _06041_ _06042_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__nor2_1
XFILLER_104_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11003_ net47 _04849_ _05143_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__a21o_1
XFILLER_93_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12954_ clknet_leaf_30_clk _00173_ VGND VGND VPWR VPWR _246_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11905_ _05888_ _05890_ _05897_ _05908_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__o31a_2
XFILLER_93_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12885_ _01233_ _01239_ _06487_ _01296_ _096_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__a32o_1
XFILLER_73_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11836_ _152_\[10\] _05844_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__or2_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11767_ _05782_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__inv_2
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13506_ clknet_leaf_60_clk _00725_ VGND VGND VPWR VPWR _152_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10718_ _173_\[13\] _04917_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__or2_1
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11698_ _05721_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10649_ _173_\[23\] _04663_ _04895_ _04891_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__o211a_1
XFILLER_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13437_ clknet_leaf_129_clk _00656_ VGND VGND VPWR VPWR _164_\[23\] sky130_fd_sc_hd__dfxtp_1
X_13368_ clknet_leaf_125_clk _00587_ VGND VGND VPWR VPWR _170_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12319_ _06191_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__clkbuf_1
X_13299_ clknet_leaf_23_clk _00518_ VGND VGND VPWR VPWR _176_\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07860_ _02342_ _02397_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__or2_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06811_ _01420_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__buf_2
X_07791_ _02327_ _02330_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__nand2_1
X_09530_ _01277_ _03878_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__nand2_4
X_06742_ net34 VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__inv_2
XFILLER_83_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09461_ _02871_ _01421_ _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06673_ _01366_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__buf_4
XFILLER_91_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09392_ _228_\[29\] _231_\[29\] _03797_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__o21a_1
X_08412_ _02852_ _01801_ _02824_ _02853_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__o211a_1
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08343_ _228_\[9\] _02775_ _02753_ _02800_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__a211o_1
XFILLER_138_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08274_ _231_\[24\] _02706_ _02695_ _02748_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__o211a_1
XFILLER_32_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07225_ _01756_ _01779_ _01785_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07156_ _01718_ _01719_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__and2_1
XFILLER_133_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07087_ _173_\[18\] _01646_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__or2_1
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09728_ _04112_ _04116_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__and2_1
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07989_ _02518_ _02523_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__and2_1
XFILLER_83_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09659_ _01278_ _01292_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__nand2_2
XFILLER_103_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12670_ _06375_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _149_\[20\] _05262_ _05652_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__a21o_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11552_ _05590_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10503_ _173_\[10\] _04780_ _04794_ _04785_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__o211a_1
X_11483_ _116_\[7\] _05527_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__nor2_1
XFILLER_7_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13222_ clknet_leaf_24_clk _00441_ VGND VGND VPWR VPWR _182_\[0\] sky130_fd_sc_hd__dfxtp_1
X_10434_ _176_\[22\] _04735_ _04745_ _04740_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__o211a_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10365_ _01216_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__buf_2
X_13153_ clknet_leaf_13_clk _00372_ VGND VGND VPWR VPWR _225_\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12104_ _06078_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__clkbuf_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10296_ _182_\[9\] _04634_ _04652_ _04649_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__o211a_1
XFILLER_97_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ clknet_leaf_100_clk _00303_ VGND VGND VPWR VPWR _234_\[28\] sky130_fd_sc_hd__dfxtp_1
X_12035_ _06010_ _06011_ _06022_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__or3_1
XFILLER_77_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13986_ clknet_leaf_31_clk _01205_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12937_ clknet_leaf_39_clk _00156_ VGND VGND VPWR VPWR _246_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12868_ _118_\[25\] _120_\[25\] _06473_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__mux2_1
XFILLER_33_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11819_ _05742_ _05829_ _05830_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__and3_1
XFILLER_61_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _122_\[24\] _120_\[24\] _06434_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__mux2_1
XFILLER_21_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07010_ _173_\[1\] _01604_ _01569_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__mux2_1
XFILLER_143_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08961_ _02833_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__buf_6
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08892_ _03290_ _03292_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__and2b_1
X_07912_ _02430_ _02431_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__and2b_1
XFILLER_111_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07843_ _01661_ _01612_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__xnor2_2
XFILLER_57_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07774_ _02314_ _02315_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__nor2_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09513_ _01235_ _03899_ _03906_ _03909_ _03910_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__o311a_1
X_06725_ _01396_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06656_ _01354_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__buf_6
X_09444_ _02871_ _231_\[31\] _228_\[31\] VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__a21o_1
XFILLER_25_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06587_ _01276_ _01292_ _01278_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09375_ _185_\[29\] _03780_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__nand2_1
X_08326_ _225_\[6\] VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__clkbuf_4
X_08257_ _164_\[19\] _02736_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__or2_1
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07208_ _01608_ _01769_ _01411_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_5_0_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_08188_ _01518_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__buf_4
XFILLER_118_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07139_ _173_\[30\] _01704_ _01672_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__mux2_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10150_ _01233_ _03903_ _03876_ _04521_ _04437_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__o311a_1
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10081_ _03901_ _04160_ _04333_ _03935_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__a211o_1
XFILLER_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13840_ clknet_leaf_95_clk _01059_ VGND VGND VPWR VPWR _126_\[16\] sky130_fd_sc_hd__dfxtp_1
X_13771_ clknet_leaf_87_clk _00990_ VGND VGND VPWR VPWR _130_\[11\] sky130_fd_sc_hd__dfxtp_1
X_10983_ net54 _04853_ _05130_ _05117_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__o211a_1
XFILLER_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12722_ _124_\[19\] _122_\[19\] _06401_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__mux2_1
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12653_ _06366_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11604_ _118_\[5\] _05636_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__xnor2_1
X_12584_ _06330_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__clkbuf_1
X_11535_ _118_\[19\] _05574_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13205_ clknet_leaf_40_clk _00424_ VGND VGND VPWR VPWR _185_\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_99_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11466_ _05511_ _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__xnor2_1
X_11397_ _149_\[28\] _132_\[28\] VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__nand2_1
X_10417_ _179_\[18\] _182_\[18\] _04693_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__mux2_1
XFILLER_140_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10348_ _04681_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__clkbuf_4
X_13136_ clknet_leaf_117_clk _00355_ VGND VGND VPWR VPWR _228_\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10279_ _179_\[3\] _04629_ _04641_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__a21o_1
XFILLER_3_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13067_ clknet_leaf_106_clk _00286_ VGND VGND VPWR VPWR _234_\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12018_ _152_\[25\] _05995_ _05996_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__nand3_1
XFILLER_78_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13969_ clknet_leaf_96_clk _01188_ VGND VGND VPWR VPWR _118_\[17\] sky130_fd_sc_hd__dfxtp_2
X_06510_ _01220_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__inv_2
XFILLER_81_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07490_ _185_\[12\] _234_\[12\] VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__or2_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09160_ _03558_ _03560_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__and2b_1
X_09091_ _03499_ _03504_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__a21oi_1
X_08111_ _02625_ _02632_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__or2_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08042_ _185_\[30\] _234_\[30\] VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__and2_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09993_ _04370_ _04371_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08944_ _03310_ _03329_ _03360_ _03361_ _03362_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__o221a_1
XFILLER_96_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08875_ _03293_ _03295_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__xor2_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07826_ _02363_ _02364_ _02362_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__a21o_1
XFILLER_72_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07757_ _182_\[20\] _01671_ _02291_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__a21o_1
X_06708_ _01386_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07688_ _01664_ _01827_ _02178_ _02232_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__a211o_1
XFILLER_40_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06639_ _01252_ _01340_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__or2_1
XFILLER_80_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09427_ _03794_ _03813_ _03831_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__o21ai_1
X_09358_ _03739_ _03740_ _03764_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__a21o_1
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08309_ _228_\[1\] _02771_ _02765_ _02774_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__o211a_1
XFILLER_126_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11320_ _05368_ _05373_ _05376_ _05383_ _05375_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__a311o_1
XFILLER_60_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09289_ _170_\[26\] _02855_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__or2_1
XFILLER_126_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11251_ _152_\[9\] _05325_ _05318_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__mux2_1
XFILLER_109_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11182_ _05263_ _05264_ _05265_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__and3_1
X_10202_ _185_\[28\] _03870_ _03864_ _04571_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__o211a_1
XFILLER_106_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10133_ _04472_ _04482_ _04504_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10064_ _01244_ _04051_ _03903_ _03952_ _03960_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__a32o_1
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13823_ clknet_leaf_65_clk _01042_ VGND VGND VPWR VPWR _128_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13754_ clknet_leaf_66_clk _00973_ VGND VGND VPWR VPWR _132_\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10966_ _164_\[21\] _05107_ _05094_ _05118_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__o211a_1
XFILLER_16_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13685_ clknet_leaf_77_clk _00904_ VGND VGND VPWR VPWR _136_\[21\] sky130_fd_sc_hd__dfxtp_1
X_10897_ net36 _05068_ _05070_ _05035_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__a211o_1
X_12705_ _124_\[11\] _122_\[11\] _06390_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__mux2_1
X_12636_ _126_\[10\] _124_\[10\] _06357_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__mux2_1
XFILLER_31_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12567_ _06321_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12498_ _06285_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__clkbuf_1
X_11518_ _05558_ _05559_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__nand2_1
XFILLER_125_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11449_ _05487_ _05490_ _05486_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__a21o_1
XFILLER_7_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13119_ clknet_leaf_119_clk _00338_ VGND VGND VPWR VPWR _231_\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06990_ _240_\[27\] _01565_ _01558_ _01590_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__o211a_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _03050_ _03052_ _03087_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__a21bo_1
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07611_ _02119_ _02121_ _02157_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__a21oi_1
XFILLER_66_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08591_ _03002_ _03003_ _03019_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07542_ _185_\[14\] _234_\[14\] VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__nand2_1
XFILLER_34_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07473_ _182_\[11\] _01638_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__or2_1
XFILLER_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09212_ _228_\[24\] _231_\[24\] _02849_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__a21o_1
X_09143_ _03519_ _03525_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__nor2_1
XFILLER_135_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09074_ _03486_ _03488_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08025_ _02557_ _02558_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__or2b_1
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09976_ _246_\[19\] _01315_ _01300_ _179_\[19\] VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__o22a_1
XFILLER_103_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08927_ _02151_ _03345_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08858_ _02858_ _03278_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__xnor2_2
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07809_ _02348_ _02349_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__nor2_2
XFILLER_45_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08789_ _03129_ _03131_ _03181_ _03182_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__a211oi_1
XFILLER_53_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10820_ _164_\[10\] _04983_ _05015_ _04998_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__o211a_1
X_10751_ _167_\[22\] _04945_ _04966_ _04952_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__a211o_1
XFILLER_13_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13470_ clknet_leaf_122_clk _00689_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfxtp_2
X_12421_ _132_\[4\] _130_\[4\] _06201_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__mux2_1
XFILLER_71_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10682_ _01216_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12352_ _06209_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__clkbuf_1
X_12283_ _06172_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__clkbuf_1
X_11303_ _05355_ _05364_ _05361_ _05360_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__a31o_1
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11234_ _152_\[7\] _05310_ _01362_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__mux2_1
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11165_ net20 _05202_ _05192_ _158_\[18\] VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__a22o_1
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11096_ _158_\[1\] _158_\[0\] _05194_ _05196_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__o31a_1
XFILLER_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10116_ _04449_ _04467_ _04489_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__a21o_1
XFILLER_95_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10047_ _04422_ _04423_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__nor2_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11998_ _142_\[24\] _05993_ _05893_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__mux2_1
XFILLER_17_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13806_ clknet_leaf_98_clk _01025_ VGND VGND VPWR VPWR _128_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13737_ clknet_leaf_58_clk _00956_ VGND VGND VPWR VPWR _132_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10949_ net43 _05068_ _05106_ _05086_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_70_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13668_ clknet_leaf_54_clk _00887_ VGND VGND VPWR VPWR _136_\[4\] sky130_fd_sc_hd__dfxtp_1
X_12619_ _126_\[2\] _124_\[2\] _06346_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__mux2_1
X_13599_ clknet_leaf_56_clk _00818_ VGND VGND VPWR VPWR _142_\[31\] sky130_fd_sc_hd__dfxtp_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09830_ _01242_ _03890_ _03896_ _03927_ _04215_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__a41o_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09761_ _185_\[9\] _03869_ _03919_ _04149_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__o211a_1
XFILLER_112_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06973_ _01568_ _01578_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__or2_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _02871_ _03137_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__xnor2_2
XFILLER_132_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09692_ _04081_ _04082_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__nor2_1
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08643_ _02835_ _02797_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ _01838_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__clkinv_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07525_ _02073_ _02074_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__xnor2_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_50_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07456_ _01661_ _01616_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07387_ _01941_ _01942_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__nor2_1
XFILLER_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09126_ _170_\[22\] _02842_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__nor2_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09057_ _03404_ _03436_ _03471_ _03462_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__and4_1
XFILLER_136_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08008_ _185_\[29\] _234_\[29\] VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__or2_1
XFILLER_2_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09959_ _04335_ _04336_ _04338_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__or3b_2
XFILLER_104_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12970_ clknet_leaf_19_clk _00189_ VGND VGND VPWR VPWR _243_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11921_ _152_\[18\] _05921_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__or2_1
XFILLER_73_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11852_ _05859_ _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__xnor2_1
X_10803_ _167_\[5\] _04980_ _04958_ _05003_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_52_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_16
X_11783_ _05796_ _05797_ net28 _05776_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__a2bb2o_1
X_13522_ clknet_leaf_80_clk _00741_ VGND VGND VPWR VPWR _152_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10734_ _170_\[17\] _04942_ _04922_ _04954_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__o211a_1
X_10665_ _04683_ _04904_ _04905_ _04891_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__o211a_1
X_13453_ clknet_leaf_2_clk _00672_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfxtp_4
X_12404_ _06236_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__clkbuf_1
X_13384_ clknet_leaf_1_clk _00603_ VGND VGND VPWR VPWR _167_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12335_ _06199_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__clkbuf_1
X_10596_ _04853_ _04858_ _04859_ _04839_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__a211o_1
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12266_ _06163_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11217_ _05289_ _05290_ _05288_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__o21ai_1
X_12197_ _06127_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11148_ _01261_ _05239_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__nand2_1
XFILLER_96_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11079_ net60 _04628_ _05189_ _05117_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__o211a_1
XFILLER_64_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_16
X_07310_ _185_\[6\] _234_\[6\] VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__nand2_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08290_ _01420_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__buf_2
X_07241_ _01437_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__buf_4
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07172_ _01733_ _01734_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09813_ _03868_ _04199_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__nand2_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09744_ _03933_ _04087_ _04132_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__or3_1
X_06956_ _240_\[17\] _01565_ _01558_ _01566_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__o211a_1
X_09675_ _04038_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__inv_2
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06887_ _243_\[30\] _01474_ _01510_ _01516_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__o211a_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _170_\[6\] _02787_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__nand2_1
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_70_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08557_ _02953_ _02955_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__nor2_1
XFILLER_23_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07508_ _02053_ _02058_ _01427_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__mux2_1
X_08488_ _01734_ _02898_ _02920_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__a21oi_1
X_07439_ _01941_ _01963_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__or2b_1
XFILLER_50_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10450_ _179_\[27\] _04721_ _04751_ _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__o211a_1
XFILLER_109_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09109_ _185_\[21\] _03521_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__or2_1
X_10381_ _176_\[7\] _04683_ _04707_ _01419_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__a211o_1
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12120_ _140_\[21\] _142_\[21\] _06079_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__mux2_1
XFILLER_2_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12051_ _06039_ _06040_ _152_\[29\] VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__a21oi_1
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11002_ _164_\[1\] net68 _02907_ _04692_ _02711_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__a221o_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12953_ clknet_leaf_21_clk _00172_ VGND VGND VPWR VPWR _246_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11904_ _152_\[15\] _05896_ _05907_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__o21ai_1
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12884_ _01276_ _01292_ _03958_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__and3_1
XFILLER_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11835_ _152_\[10\] _05844_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__nand2_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_60_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11766_ _05780_ _05781_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__nand2_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13505_ clknet_leaf_57_clk _00724_ VGND VGND VPWR VPWR _152_\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ _01225_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__buf_2
X_11697_ _149_\[28\] _05720_ _05625_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__mux2_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13436_ clknet_leaf_122_clk _00655_ VGND VGND VPWR VPWR _164_\[22\] sky130_fd_sc_hd__dfxtp_1
X_10648_ _02359_ _04894_ _04630_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__mux2_1
X_10579_ _04637_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__buf_4
X_13367_ clknet_leaf_125_clk _00586_ VGND VGND VPWR VPWR _170_\[17\] sky130_fd_sc_hd__dfxtp_1
X_12318_ _136_\[19\] _134_\[19\] _06189_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__mux2_1
X_13298_ clknet_leaf_26_clk _00517_ VGND VGND VPWR VPWR _176_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12249_ _06154_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06810_ _01435_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__buf_2
X_07790_ _02327_ _02330_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__or2_1
X_06741_ net34 VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__inv_2
XFILLER_49_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09460_ _01423_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__buf_6
X_06672_ _01272_ _01274_ _01359_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__and3_2
XFILLER_52_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08411_ net53 _01519_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__or2_1
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09391_ _228_\[29\] _231_\[29\] _02865_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__a21o_1
XFILLER_17_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08342_ _02797_ _02791_ _02760_ _02799_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__o211a_1
X_08273_ _02686_ _02747_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__or2_1
XFILLER_20_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07224_ _01781_ _01784_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__xor2_1
XFILLER_20_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07155_ _243_\[0\] _240_\[0\] _237_\[0\] VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__mux2_1
XFILLER_145_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07086_ _237_\[18\] VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__clkbuf_8
XFILLER_121_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07988_ _02402_ _02466_ _02519_ _02522_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__o31a_1
X_09727_ _04112_ _04116_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__nor2_1
XFILLER_87_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06939_ _243_\[12\] _01536_ _01509_ _01554_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__a211o_1
XFILLER_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09658_ _03957_ _03887_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__nand2_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09589_ _01283_ _03983_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__nand2_4
X_08609_ _185_\[5\] _03006_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__nand2_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11620_ _01362_ _05650_ _05651_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__and3_1
XFILLER_70_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11551_ _149_\[13\] _05589_ _05533_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__mux2_1
XFILLER_11_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10502_ _04766_ _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__or2_1
XFILLER_11_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11482_ _118_\[10\] _05526_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13221_ clknet_leaf_38_clk _00440_ VGND VGND VPWR VPWR _185_\[31\] sky130_fd_sc_hd__dfxtp_2
XFILLER_109_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10433_ _04712_ _04744_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__or2_1
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10364_ _176_\[2\] _04691_ _04695_ _04677_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__o211a_1
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13152_ clknet_leaf_116_clk _00371_ VGND VGND VPWR VPWR _225_\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12103_ _140_\[13\] _142_\[13\] _06068_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__mux2_1
XFILLER_124_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10295_ _179_\[9\] _04646_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__or2_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ clknet_leaf_107_clk _00302_ VGND VGND VPWR VPWR _234_\[27\] sky130_fd_sc_hd__dfxtp_1
X_12034_ _06026_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13985_ clknet_leaf_31_clk _01204_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12936_ clknet_leaf_40_clk _00155_ VGND VGND VPWR VPWR _246_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12867_ _06478_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__clkbuf_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _05825_ _05828_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__or2_1
XFILLER_33_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12798_ _06442_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__clkbuf_1
X_11749_ _05766_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13419_ clknet_leaf_12_clk _00638_ VGND VGND VPWR VPWR _164_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
X_08960_ _02820_ _03032_ _03309_ _03378_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__a211o_1
X_08891_ _03296_ _03299_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__or2_1
X_07911_ _01421_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07842_ _02370_ _02371_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__and2b_1
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09512_ _195_\[5\] VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__inv_2
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07773_ _02268_ _02301_ _02312_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__nor3_1
XFILLER_37_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06724_ _118_\[25\] _116_\[25\] _01394_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__mux2_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06655_ _01353_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__buf_6
XFILLER_80_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09443_ _02807_ _02772_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__xnor2_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09374_ _02871_ _03779_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06586_ _01291_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__clkbuf_4
X_08325_ _228_\[5\] _02771_ _02765_ _02786_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__o211a_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08256_ _01339_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__buf_2
XFILLER_20_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07207_ _01751_ _01768_ _01518_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__mux2_1
XFILLER_4_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08187_ _01405_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__buf_2
XFILLER_118_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07138_ _237_\[30\] VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__buf_6
XFILLER_145_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07069_ _173_\[14\] _01646_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__or2_1
XFILLER_0_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10080_ _185_\[22\] _03870_ _03864_ _04455_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__o211a_1
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13770_ clknet_leaf_87_clk _00989_ VGND VGND VPWR VPWR _130_\[10\] sky130_fd_sc_hd__dfxtp_1
X_10982_ _05079_ _05129_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__or2_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12721_ _06402_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__clkbuf_1
X_12652_ _126_\[18\] _124_\[18\] _06357_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__mux2_1
X_11603_ _118_\[22\] _118_\[26\] VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12583_ _128_\[17\] _126_\[17\] _06324_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__mux2_1
X_11534_ _118_\[15\] _118_\[30\] VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11465_ _05501_ _05506_ _05504_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__o21ai_1
XFILLER_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13204_ clknet_leaf_36_clk _00423_ VGND VGND VPWR VPWR _185_\[14\] sky130_fd_sc_hd__dfxtp_2
X_10416_ _176_\[17\] _04725_ _04732_ _04728_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__a211o_1
X_11396_ _05444_ _05449_ _05450_ _05451_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__or4_1
XFILLER_98_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10347_ _04635_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__buf_4
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13135_ clknet_leaf_117_clk _00354_ VGND VGND VPWR VPWR _228_\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10278_ _182_\[3\] _01218_ _04631_ _03309_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__a31o_1
X_13066_ clknet_leaf_110_clk _00285_ VGND VGND VPWR VPWR _234_\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12017_ _05986_ _05999_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__or2_1
XFILLER_120_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13968_ clknet_leaf_96_clk _01187_ VGND VGND VPWR VPWR _118_\[16\] sky130_fd_sc_hd__dfxtp_4
X_12919_ clknet_leaf_73_clk _00143_ VGND VGND VPWR VPWR _116_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13899_ clknet_leaf_95_clk _01118_ VGND VGND VPWR VPWR _122_\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09090_ _03499_ _03504_ _01523_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__o21ai_1
X_08110_ _167_\[9\] _231_\[9\] _02626_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__mux2_1
XFILLER_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08041_ _185_\[30\] _234_\[30\] VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__nor2_1
XFILLER_134_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09992_ _142_\[18\] _04340_ _04341_ _04339_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08943_ _03330_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_15_0_clk clknet_3_7_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_130_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08874_ _03260_ _03262_ _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__o21a_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07825_ _02362_ _02363_ _02364_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__nand3_1
XFILLER_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07756_ _02296_ _02297_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__nand2_2
XFILLER_84_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06707_ _118_\[18\] _116_\[18\] _01381_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__mux2_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07687_ _01801_ _02224_ _02231_ _02202_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__o211a_1
XFILLER_44_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09426_ _03829_ _03830_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__nor2_1
X_06638_ _01297_ _01339_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__nor2_1
X_06569_ _01277_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__clkbuf_4
XFILLER_100_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09357_ _03762_ _03763_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__nand2_1
XFILLER_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08308_ _02749_ _02773_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__or2_1
X_09288_ _03691_ _03695_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__or2_1
XFILLER_138_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08239_ _164_\[14\] _02701_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__or2_1
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11250_ _05322_ _05324_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11181_ _149_\[0\] _132_\[0\] VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__or2_1
X_10201_ _04568_ _04570_ _03868_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__o21ai_1
XFILLER_109_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10132_ _04472_ _04482_ _04504_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__o21bai_1
XFILLER_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10063_ _04059_ _04438_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__nand2_1
XFILLER_88_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13822_ clknet_leaf_69_clk _01041_ VGND VGND VPWR VPWR _128_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13753_ clknet_leaf_67_clk _00972_ VGND VGND VPWR VPWR _132_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12704_ _06393_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__clkbuf_1
X_10965_ _167_\[21\] _05089_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__or2_1
X_13684_ clknet_leaf_77_clk _00903_ VGND VGND VPWR VPWR _136_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10896_ _164_\[0\] _05059_ _05043_ _05069_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__o211a_1
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12635_ _01392_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__buf_4
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12566_ _128_\[9\] _126_\[9\] _06313_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__mux2_1
XFILLER_129_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11517_ _116_\[10\] _05557_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__or2_1
X_12497_ _130_\[8\] _128_\[8\] _06280_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__mux2_1
XFILLER_116_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11448_ _05495_ _05496_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__or2b_1
XFILLER_124_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11379_ _05429_ _05436_ _05427_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__o21a_1
XFILLER_140_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13118_ clknet_leaf_103_clk _00337_ VGND VGND VPWR VPWR _231_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13049_ clknet_leaf_85_clk _00268_ VGND VGND VPWR VPWR _237_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08590_ _03002_ _03003_ _03019_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__nor3_1
X_07610_ _02155_ _02156_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__nand2_1
XFILLER_26_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07541_ _185_\[14\] _234_\[14\] VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__or2_1
Xclkbuf_3_4_0_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_19_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07472_ _182_\[11\] _01638_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__nand2_1
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09211_ _03620_ _03621_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__xor2_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09142_ _02337_ _03554_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09073_ _02242_ _03445_ _03487_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__o21ai_1
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08024_ _182_\[29\] _01701_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__nand2_1
XFILLER_116_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09975_ _243_\[19\] _04129_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__or2_1
XFILLER_97_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08926_ _185_\[16\] _03344_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08857_ _02820_ _02781_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__xnor2_1
X_07808_ _182_\[22\] _01678_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__and2_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08788_ _03210_ _03211_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__or2_1
X_07739_ _02275_ _02281_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__xor2_1
XFILLER_41_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10750_ _170_\[22\] _04942_ _04958_ _04965_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__o211a_1
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09409_ _02573_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__inv_2
X_10681_ _167_\[2\] _04818_ _04916_ _04891_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__o211a_1
X_12420_ _06244_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12351_ _132_\[2\] _134_\[2\] _06208_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__mux2_1
XFILLER_5_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12282_ _136_\[2\] _134_\[2\] _06167_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__mux2_1
XFILLER_138_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11302_ _05368_ _05369_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__nand2_1
XFILLER_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11233_ _05308_ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11164_ _01264_ _05251_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__nand2_1
X_11095_ net2 _05196_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__nor2_1
X_10115_ _04447_ _04465_ _04466_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__o21bai_2
XFILLER_48_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10046_ _04413_ _04421_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__and2_1
XFILLER_0_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11997_ net17 _05992_ _05785_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__mux2_1
XFILLER_90_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13805_ clknet_leaf_93_clk _01024_ VGND VGND VPWR VPWR _128_\[13\] sky130_fd_sc_hd__dfxtp_1
X_13736_ clknet_leaf_55_clk _00955_ VGND VGND VPWR VPWR _132_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10948_ _164_\[16\] _05059_ _05094_ _05105_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__o211a_1
XFILLER_31_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13667_ clknet_leaf_59_clk _00886_ VGND VGND VPWR VPWR _136_\[3\] sky130_fd_sc_hd__dfxtp_1
X_10879_ _170_\[28\] _05036_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__or2_1
X_13598_ clknet_leaf_51_clk _00817_ VGND VGND VPWR VPWR _142_\[30\] sky130_fd_sc_hd__dfxtp_1
X_12618_ _06348_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12549_ _128_\[1\] _126_\[1\] _06302_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__mux2_1
XFILLER_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 _01274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _03868_ _04148_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__nand2_1
XFILLER_58_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06972_ _176_\[22\] _240_\[22\] _01569_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__mux2_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _01278_ _03878_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__nor2_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _02842_ _02804_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08642_ _03044_ _03045_ _03046_ _03043_ _03041_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__o32ai_4
XFILLER_54_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08573_ _02990_ _02992_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__and2b_1
XFILLER_42_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07524_ _243_\[13\] _240_\[13\] _01645_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__mux2_2
XFILLER_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07455_ _02006_ _01980_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__or2_1
X_07386_ _01901_ _01926_ _01940_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__nor3_1
X_09125_ _02839_ _01426_ _03379_ _03538_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__o211a_1
X_09056_ _03371_ _03403_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__nand2_1
XFILLER_123_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08007_ _185_\[29\] _234_\[29\] VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__nand2_1
XFILLER_144_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09958_ _01284_ _04321_ _04161_ _04337_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__a211o_1
XFILLER_66_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08909_ _03288_ _03312_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__nor3_1
X_09889_ _04271_ _04272_ _03946_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__a21o_1
XFILLER_85_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11920_ _152_\[18\] _05921_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__nand2_1
XFILLER_73_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11851_ _05836_ _05847_ _05849_ _05845_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__o31ai_2
XFILLER_73_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11782_ _05780_ _05786_ _05795_ _01274_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__a31o_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10802_ _170_\[5\] _05002_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__or2_1
XFILLER_26_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13521_ clknet_leaf_81_clk _00740_ VGND VGND VPWR VPWR _152_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10733_ _173_\[17\] _04953_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__or2_1
XFILLER_41_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13452_ clknet_leaf_113_clk _00671_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfxtp_2
X_10664_ _02561_ _04724_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__nand2_1
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12403_ _132_\[27\] _134_\[27\] _06230_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__mux2_1
X_10595_ _01863_ _04631_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__nor2_1
X_13383_ clknet_leaf_12_clk _00602_ VGND VGND VPWR VPWR _167_\[1\] sky130_fd_sc_hd__dfxtp_1
X_12334_ _136_\[27\] _134_\[27\] _06189_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__mux2_1
XFILLER_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12265_ _138_\[26\] _136_\[26\] _06156_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__mux2_1
XFILLER_99_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11216_ _05293_ _05294_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__nand2_1
X_12196_ _140_\[25\] _138_\[25\] _06123_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__mux2_1
Xoutput60 net60 VGND VGND VPWR VPWR dout[31] sky130_fd_sc_hd__buf_2
X_11147_ _158_\[13\] _01260_ _158_\[14\] VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11078_ _03862_ _04724_ _05188_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__a21o_1
X_10029_ _04395_ _04405_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__nand2_1
XFILLER_48_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13719_ clknet_leaf_67_clk _00938_ VGND VGND VPWR VPWR _134_\[23\] sky130_fd_sc_hd__dfxtp_1
X_07240_ _01612_ _01649_ _01693_ _01800_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__a211o_1
X_07171_ _243_\[1\] _240_\[1\] _01604_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__mux2_2
XFILLER_145_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09812_ _04196_ _04198_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__xor2_1
XFILLER_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09743_ _03961_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__clkbuf_4
X_06955_ _176_\[17\] _01531_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__or2_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09674_ _04065_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__inv_2
X_06886_ _179_\[30\] _01302_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__or2_1
XFILLER_55_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08625_ _170_\[6\] _02787_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__or2_1
XFILLER_82_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _01814_ _02986_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07507_ _02056_ _02057_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__or2_2
XFILLER_54_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08487_ _02894_ _02897_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__nor2_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07438_ _01989_ _01990_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__nand2_1
XFILLER_136_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07369_ _01864_ _01879_ _01880_ _01911_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__and4_1
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09108_ _185_\[21\] _03521_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__nand2_1
XFILLER_108_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10380_ _179_\[7\] _04684_ _04705_ _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__o211a_1
XFILLER_123_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09039_ _228_\[19\] _231_\[19\] _03454_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__o21a_1
X_12050_ _152_\[29\] _06039_ _06040_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__and3_1
XFILLER_132_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11001_ _04855_ _05141_ _05142_ _05122_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__a211o_1
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12952_ clknet_leaf_21_clk _00171_ VGND VGND VPWR VPWR _246_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11903_ _152_\[14\] _05885_ _05896_ _152_\[15\] VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__a22o_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12883_ net25 _05196_ _06486_ _01425_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__o211a_1
XFILLER_61_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11834_ _140_\[20\] _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__xnor2_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11765_ _152_\[4\] _05779_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__or2_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13504_ clknet_leaf_56_clk _00723_ VGND VGND VPWR VPWR _152_\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _05715_ _05719_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__xor2_1
XFILLER_41_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10716_ _167_\[12\] _04836_ _04941_ _04914_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__a211o_1
XFILLER_139_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10647_ _176_\[23\] _01216_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__or2_1
X_13435_ clknet_leaf_125_clk _00654_ VGND VGND VPWR VPWR _164_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10578_ _04691_ _04846_ _04847_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__a21o_1
X_13366_ clknet_leaf_125_clk _00585_ VGND VGND VPWR VPWR _170_\[16\] sky130_fd_sc_hd__dfxtp_1
X_12317_ _06190_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__clkbuf_1
X_13297_ clknet_leaf_24_clk _00516_ VGND VGND VPWR VPWR _176_\[11\] sky130_fd_sc_hd__dfxtp_1
X_12248_ _138_\[18\] _136_\[18\] _06145_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__mux2_1
XFILLER_122_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12179_ _140_\[17\] _138_\[17\] _06112_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__mux2_1
XFILLER_96_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06740_ net34 VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__inv_2
XFILLER_110_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06671_ _01365_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08410_ _225_\[25\] VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__buf_4
XFILLER_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09390_ _03794_ _03795_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__or2_1
XFILLER_36_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08341_ net67 _02798_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__or2_1
X_08272_ _164_\[24\] _228_\[24\] _02687_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__mux2_1
XFILLER_20_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07223_ _01782_ _01783_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__nand2_1
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07154_ _01714_ _01717_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07085_ _240_\[17\] _01660_ _01653_ _01663_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__o211a_1
XFILLER_133_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07987_ _02463_ _02497_ _02519_ _02520_ _02521_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__o221a_1
XFILLER_47_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09726_ _04114_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__or2_1
XFILLER_86_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06938_ _240_\[12\] _01526_ _01510_ _01553_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__o211a_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09657_ _04047_ _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__or2_1
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06869_ _243_\[25\] _01474_ _01461_ _01503_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__o211a_1
XFILLER_70_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09588_ _01279_ _03874_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__nor2b_4
X_08608_ _03033_ _03036_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__xnor2_2
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _01856_ _02946_ _02970_ _02355_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__a211o_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11550_ _05587_ _05588_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10501_ _176_\[10\] _179_\[10\] _04790_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__mux2_1
XFILLER_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13220_ clknet_leaf_37_clk _00439_ VGND VGND VPWR VPWR _185_\[30\] sky130_fd_sc_hd__dfxtp_2
X_11481_ _118_\[25\] _118_\[14\] VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10432_ _179_\[22\] _182_\[22\] _04743_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__mux2_1
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10363_ _04692_ _04694_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__or2_1
X_13151_ clknet_leaf_104_clk _00370_ VGND VGND VPWR VPWR _228_\[31\] sky130_fd_sc_hd__dfxtp_1
X_12102_ _06077_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13082_ clknet_leaf_102_clk _00301_ VGND VGND VPWR VPWR _234_\[26\] sky130_fd_sc_hd__dfxtp_1
X_12033_ _142_\[27\] _06025_ _06005_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__mux2_1
X_10294_ _179_\[8\] _04629_ _04651_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__a21o_1
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13984_ clknet_leaf_36_clk _01203_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12935_ clknet_leaf_40_clk _00154_ VGND VGND VPWR VPWR _246_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _118_\[24\] _120_\[24\] _06473_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__mux2_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _05825_ _05828_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__nand2_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _122_\[23\] _120_\[23\] _06434_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__mux2_1
X_11748_ _142_\[2\] _05764_ _05765_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__mux2_1
XFILLER_14_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11679_ _118_\[13\] _05703_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__xnor2_1
X_13418_ clknet_leaf_3_clk _00637_ VGND VGND VPWR VPWR _164_\[4\] sky130_fd_sc_hd__dfxtp_1
X_13349_ clknet_leaf_8_clk _00568_ VGND VGND VPWR VPWR _173_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07910_ _01687_ _01973_ _02419_ _02447_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__o211a_1
X_08890_ _03295_ _03293_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__or2b_1
XFILLER_69_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07841_ _01437_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__buf_4
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07772_ _02313_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__inv_2
X_09511_ _03880_ _03908_ _01235_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__o21ai_1
XFILLER_110_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06723_ _01395_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06654_ _01302_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__buf_4
XFILLER_80_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09442_ _02582_ _03823_ _03821_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__a21oi_1
X_06585_ _195_\[1\] _195_\[0\] VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__and2_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09373_ _02830_ _02801_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08324_ _02749_ _02785_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__or2_1
XFILLER_33_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08255_ _231_\[18\] _02730_ _02712_ _02735_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__a211o_1
XFILLER_137_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07206_ _01766_ _01767_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__nor2_1
X_08186_ _234_\[31\] _02646_ _02664_ _02685_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__a211o_1
XFILLER_133_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07137_ _240_\[29\] _01660_ _01653_ _01703_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__o211a_1
XFILLER_4_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07068_ _237_\[14\] VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__buf_4
XFILLER_133_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09709_ _185_\[7\] _03869_ _03919_ _04099_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__o211a_1
XFILLER_83_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10981_ _164_\[26\] _167_\[26\] _01214_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__mux2_1
XFILLER_74_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12720_ _124_\[18\] _122_\[18\] _06401_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__mux2_1
XFILLER_130_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12651_ _06365_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11602_ _149_\[18\] _05352_ _05634_ _05635_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__a22o_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12582_ _06329_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__clkbuf_1
X_11533_ _05573_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11464_ _116_\[5\] _05510_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13203_ clknet_leaf_36_clk _00422_ VGND VGND VPWR VPWR _185_\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_99_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10415_ _179_\[17\] _04721_ _04705_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__o211a_1
X_11395_ _05443_ _05434_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__and2b_1
X_10346_ _182_\[31\] _04663_ _04680_ _04677_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__o211a_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13134_ clknet_leaf_115_clk _00353_ VGND VGND VPWR VPWR _228_\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10277_ _182_\[2\] _04634_ _04640_ _00105_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__o211a_1
X_13065_ clknet_leaf_109_clk _00284_ VGND VGND VPWR VPWR _234_\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12016_ _06008_ _06009_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__nand2_1
XFILLER_39_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13967_ clknet_leaf_97_clk _01186_ VGND VGND VPWR VPWR _118_\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_74_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12918_ clknet_leaf_87_clk _00142_ VGND VGND VPWR VPWR _116_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13898_ clknet_leaf_97_clk _01117_ VGND VGND VPWR VPWR _122_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12849_ _118_\[16\] _120_\[16\] _06462_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__mux2_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08040_ _01681_ _02572_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__xnor2_4
XFILLER_128_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09991_ _04358_ _04369_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08942_ _03251_ _03297_ _03298_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__a21o_1
XFILLER_130_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08873_ _03263_ _03265_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__or2b_1
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07824_ _185_\[23\] _234_\[23\] VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__nand2_1
X_07755_ _182_\[21\] _01675_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__or2_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07686_ _01409_ _02230_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__nand2_1
X_06706_ _01385_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06637_ _01302_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__buf_4
XFILLER_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09425_ _03825_ _03826_ _03828_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__a21oi_1
XFILLER_13_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06568_ _195_\[2\] VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__buf_2
X_09356_ _03722_ _03741_ _03761_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__or3_1
X_06499_ _01212_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__inv_2
XFILLER_100_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08307_ net47 _02772_ _02750_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__mux2_1
X_09287_ _03691_ _03695_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__nand2_1
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08238_ _01420_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__clkbuf_4
XFILLER_118_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10200_ _04567_ _04569_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__and2_1
X_08169_ _231_\[26\] _02649_ _02641_ _02673_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__o211a_1
XFILLER_134_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11180_ _149_\[0\] _132_\[0\] VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__nand2_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10131_ _04497_ _04503_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10062_ _04436_ _04160_ _04437_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__a21oi_1
XFILLER_121_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13821_ clknet_leaf_68_clk _01040_ VGND VGND VPWR VPWR _128_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13752_ clknet_leaf_67_clk _00971_ VGND VGND VPWR VPWR _132_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10964_ net48 _04853_ _05116_ _05117_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__o211a_1
X_12703_ _124_\[10\] _122_\[10\] _06390_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__mux2_1
X_13683_ clknet_leaf_77_clk _00902_ VGND VGND VPWR VPWR _136_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10895_ _167_\[0\] _05036_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__or2_1
X_12634_ _06356_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__clkbuf_1
X_12565_ _06320_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11516_ _116_\[10\] _05557_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__nand2_1
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12496_ _06284_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11447_ _116_\[3\] _05494_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__or2_1
XFILLER_125_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11378_ _149_\[24\] _132_\[24\] _149_\[25\] _132_\[25\] VGND VGND VPWR VPWR _05436_
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10329_ _179_\[24\] _04658_ _04670_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__a21o_1
X_13117_ clknet_leaf_119_clk _00336_ VGND VGND VPWR VPWR _231_\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13048_ clknet_leaf_110_clk _00267_ VGND VGND VPWR VPWR _237_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07540_ _01687_ _02088_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07471_ _01989_ _01994_ _02021_ _01923_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__a31o_1
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09210_ _02371_ _03580_ _03578_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__a21bo_1
X_09141_ _03552_ _03553_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__xnor2_1
X_09072_ _185_\[19\] _03444_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__nand2_1
XFILLER_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08023_ _182_\[29\] _01701_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__nor2_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09974_ _185_\[18\] _04150_ _04175_ _04353_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__o211a_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08925_ _02865_ _03343_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08856_ _02811_ _03032_ _02861_ _03277_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__a211o_1
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07807_ _182_\[22\] _01678_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__nor2_1
XFILLER_45_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08787_ _170_\[11\] _02804_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__nor2_1
X_07738_ _02148_ _02278_ _02280_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__a21bo_1
XFILLER_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07669_ _02186_ _02206_ _02212_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__and3_1
XFILLER_80_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09408_ _03796_ _03798_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__and2b_1
XFILLER_25_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10680_ _04888_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__or2_1
XFILLER_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09339_ _185_\[28\] _03745_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__nand2_1
XFILLER_139_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12350_ _06004_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__buf_4
XFILLER_5_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12281_ _06171_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11301_ _149_\[16\] _132_\[16\] VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__or2_1
X_11232_ _05301_ _05303_ _05300_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__o21ai_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11163_ _158_\[18\] _01263_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__nand2_1
XFILLER_106_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10114_ _04486_ _04487_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__nor2_1
XFILLER_96_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11094_ _158_\[1\] VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__inv_2
XFILLER_121_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10045_ _04413_ _04421_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__nor2_1
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13804_ clknet_leaf_87_clk _01023_ VGND VGND VPWR VPWR _128_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11996_ _05986_ _05991_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__xor2_1
XFILLER_91_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13735_ clknet_leaf_59_clk _00954_ VGND VGND VPWR VPWR _132_\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10947_ _167_\[16\] _05089_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__or2_1
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13666_ clknet_leaf_54_clk _00885_ VGND VGND VPWR VPWR _136_\[2\] sky130_fd_sc_hd__dfxtp_1
X_12617_ _126_\[1\] _124_\[1\] _06346_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__mux2_1
X_10878_ _164_\[27\] _05025_ _05056_ _05035_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__a211o_1
X_13597_ clknet_leaf_36_clk _00816_ VGND VGND VPWR VPWR _142_\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_14_0_clk clknet_3_7_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_129_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12548_ _06311_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12479_ _06275_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 _01302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06971_ _243_\[21\] _01548_ _01545_ _01577_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__o211a_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _03884_ _03898_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__nand2_1
X_08710_ _03111_ _03112_ _03113_ _03110_ _03109_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__o32ai_4
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08641_ _03068_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__inv_2
XFILLER_27_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08572_ _02987_ _02989_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__nor2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07523_ _02070_ _02072_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07454_ _01977_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__inv_2
XFILLER_62_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07385_ _01901_ _01926_ _01940_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__o21a_1
XFILLER_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09124_ _01428_ _03512_ _03537_ _01495_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__a211o_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09055_ _03372_ _03405_ _03436_ _03462_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__or4bb_1
X_08006_ _01678_ _02539_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__xnor2_4
XFILLER_144_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09957_ _01243_ _03897_ _04005_ _03925_ _04051_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__o311a_1
XFILLER_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08908_ _03325_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__xnor2_1
X_09888_ _04266_ _04270_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__or2_1
XFILLER_106_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08839_ _03223_ _03225_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__nor2_1
XFILLER_58_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11850_ _05857_ _05858_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__or2b_1
XFILLER_122_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11781_ _05780_ _05786_ _05795_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__a21oi_1
XFILLER_82_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10801_ _01216_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__clkbuf_2
X_13520_ clknet_leaf_79_clk _00739_ VGND VGND VPWR VPWR _152_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10732_ _01216_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__clkbuf_2
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13451_ clknet_leaf_12_clk _00670_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfxtp_4
XFILLER_41_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10663_ _173_\[29\] _176_\[29\] _01226_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__mux2_1
XFILLER_13_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12402_ _06235_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__clkbuf_1
X_10594_ _173_\[6\] _176_\[6\] _01226_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__mux2_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13382_ clknet_leaf_0_clk _00601_ VGND VGND VPWR VPWR _167_\[0\] sky130_fd_sc_hd__dfxtp_1
X_12333_ _06198_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_5_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12264_ _06162_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput50 net50 VGND VGND VPWR VPWR dout[22] sky130_fd_sc_hd__buf_2
X_11215_ _149_\[5\] _132_\[5\] VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__nand2_1
X_12195_ _06126_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput61 net61 VGND VGND VPWR VPWR dout[3] sky130_fd_sc_hd__buf_2
X_11146_ _05227_ _05237_ _05238_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__a21o_1
XFILLER_68_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11077_ _164_\[31\] _01217_ _04630_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__o21a_1
X_10028_ _04395_ _04405_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__or2_1
XFILLER_49_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13718_ clknet_leaf_67_clk _00937_ VGND VGND VPWR VPWR _134_\[22\] sky130_fd_sc_hd__dfxtp_1
X_11979_ _05974_ _05975_ _152_\[23\] VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13649_ clknet_leaf_78_clk _00868_ VGND VGND VPWR VPWR _138_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07170_ _01731_ _01732_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_120_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_120_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_145_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09811_ _04144_ _04151_ _04171_ _04197_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__a31o_1
XFILLER_87_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09742_ _142_\[9\] _04130_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06954_ _01427_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__buf_2
X_09673_ _04063_ _04064_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__xnor2_1
X_06885_ _246_\[29\] _01485_ _01481_ _01515_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__o211a_1
XFILLER_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08624_ _03050_ _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__xor2_1
XFILLER_70_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _02983_ _02985_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07506_ _02055_ _02054_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__and2b_1
X_08486_ _01762_ _02918_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07437_ _01986_ _01988_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__or2_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07368_ _01877_ _01908_ _01909_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__o21a_1
XFILLER_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09107_ _02846_ _03520_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07299_ _182_\[6\] _01623_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_111_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_111_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09038_ _228_\[19\] _231_\[19\] _02830_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__a21o_1
XFILLER_89_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11000_ _02886_ _04631_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__nor2_1
XFILLER_132_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12951_ clknet_leaf_22_clk _00170_ VGND VGND VPWR VPWR _246_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12882_ _099_ _05190_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__or2_1
X_11902_ _05904_ _05905_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__nand2_1
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11833_ _140_\[27\] _140_\[29\] VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__xnor2_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _152_\[4\] _05779_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__nand2_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13503_ clknet_leaf_37_clk _00722_ VGND VGND VPWR VPWR _158_\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _05683_ _05697_ _05716_ _05718_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__o31a_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10715_ _170_\[12\] _04833_ _04922_ _04940_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__o211a_1
X_10646_ _173_\[22\] _04663_ _04893_ _04891_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__o211a_1
X_13434_ clknet_leaf_130_clk _00653_ VGND VGND VPWR VPWR _164_\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10577_ _01711_ _01712_ _04724_ _01710_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_102_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_102_clk sky130_fd_sc_hd__clkbuf_16
X_13365_ clknet_leaf_124_clk _00584_ VGND VGND VPWR VPWR _170_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12316_ _136_\[18\] _134_\[18\] _06189_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__mux2_1
X_13296_ clknet_leaf_26_clk _00515_ VGND VGND VPWR VPWR _176_\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12247_ _06153_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12178_ _06117_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__clkbuf_1
X_11129_ _05224_ _05225_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__or2_1
XFILLER_84_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06670_ _116_\[2\] _118_\[2\] _01362_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__mux2_1
XFILLER_91_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08340_ _01339_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__clkbuf_2
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08271_ _231_\[23\] _02706_ _02695_ _02746_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__o211a_1
X_07222_ _185_\[3\] _234_\[3\] VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__or2_1
XFILLER_118_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07153_ _01715_ _01716_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__nand2_1
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07084_ _01615_ _01662_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__or2_1
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07986_ _02498_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__inv_2
X_09725_ _142_\[8\] _04113_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__nor2_1
XFILLER_101_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06937_ _176_\[12\] _01531_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__or2_1
XFILLER_28_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09656_ _04045_ _04046_ _142_\[6\] VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__a21oi_1
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06868_ _179_\[25\] _01301_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__or2_1
X_08607_ _185_\[6\] _03035_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09587_ _01240_ _01278_ _01291_ _01234_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__o31a_1
X_06799_ _179_\[7\] _01300_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__or2_1
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _01923_ _02968_ _02969_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__nor3_1
X_08469_ _02900_ _02902_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__xor2_1
XFILLER_23_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10500_ _173_\[9\] _04780_ _04792_ _04785_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__o211a_1
XFILLER_137_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11480_ _05525_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10431_ _01214_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__buf_4
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10362_ _179_\[2\] _182_\[2\] _04693_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__mux2_1
X_13150_ clknet_leaf_120_clk _00369_ VGND VGND VPWR VPWR _228_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12101_ _140_\[12\] _142_\[12\] _06068_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__mux2_1
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10293_ _182_\[8\] _01218_ _04642_ _04650_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__a31o_1
XFILLER_88_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13081_ clknet_leaf_99_clk _00300_ VGND VGND VPWR VPWR _234_\[25\] sky130_fd_sc_hd__dfxtp_1
X_12032_ net20 _06024_ _05785_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__mux2_1
XFILLER_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13983_ clknet_leaf_68_clk _01202_ VGND VGND VPWR VPWR _118_\[31\] sky130_fd_sc_hd__dfxtp_2
XFILLER_19_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12934_ clknet_leaf_39_clk _00153_ VGND VGND VPWR VPWR _246_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12865_ _06477_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _05815_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__or2_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _06441_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__clkbuf_1
X_11747_ _01361_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__clkbuf_4
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11678_ _118_\[30\] _118_\[2\] VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10629_ _02181_ _04724_ _04848_ _173_\[17\] _04881_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__a221o_1
X_13417_ clknet_leaf_1_clk _00636_ VGND VGND VPWR VPWR _164_\[3\] sky130_fd_sc_hd__dfxtp_1
X_13348_ clknet_leaf_11_clk _00567_ VGND VGND VPWR VPWR _173_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13279_ clknet_leaf_7_clk _00498_ VGND VGND VPWR VPWR _179_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07840_ _01681_ _01973_ _01886_ _02379_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__o211a_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07771_ _02268_ _02301_ _02312_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__o21ai_1
X_09510_ _01283_ _03907_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__nor2_1
XFILLER_77_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06722_ _118_\[24\] _116_\[24\] _01394_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__mux2_1
X_06653_ _01303_ _01342_ _01340_ _01352_ VGND VGND VPWR VPWR _436_\[3\] sky130_fd_sc_hd__a211o_1
XFILLER_52_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09441_ _03826_ _03828_ _03825_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__a21bo_1
XFILLER_24_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06584_ _01286_ _01290_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__nor2_1
XFILLER_91_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09372_ _02506_ _03746_ _03747_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__nand3_1
XFILLER_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08323_ net63 _02784_ _02750_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__mux2_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08254_ _228_\[18\] _02733_ _02723_ _02734_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__o211a_1
XFILLER_119_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07205_ _01764_ _01765_ _01736_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__a21oi_1
X_08185_ _231_\[31\] _02649_ _02679_ _02684_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__o211a_1
XFILLER_134_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07136_ _01670_ _01702_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__or2_1
X_07067_ _01495_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__clkbuf_4
XFILLER_133_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09708_ _04095_ _04097_ _04098_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__a21o_1
XFILLER_114_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07969_ _02494_ _02495_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__and2b_1
XFILLER_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10980_ net53 _05110_ _05128_ _05122_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__a211o_1
X_09639_ _03977_ _04031_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__nor2_1
XFILLER_83_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12650_ _126_\[17\] _124_\[17\] _06357_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__mux2_1
X_11601_ _05631_ _05633_ _05352_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12581_ _128_\[16\] _126_\[16\] _06324_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__mux2_1
XFILLER_129_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11532_ _149_\[11\] _05572_ _05533_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__mux2_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11463_ _118_\[8\] _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13202_ clknet_leaf_35_clk _00421_ VGND VGND VPWR VPWR _185_\[12\] sky130_fd_sc_hd__dfxtp_2
X_10414_ _182_\[17\] _04696_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__or2_1
XFILLER_136_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11394_ _05427_ _05441_ _05436_ _05445_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__and4_1
XFILLER_99_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13133_ clknet_leaf_117_clk _00352_ VGND VGND VPWR VPWR _228_\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10345_ _179_\[31\] _04637_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__or2_1
XFILLER_140_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10276_ _179_\[2\] _04638_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__or2_1
XFILLER_97_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13064_ clknet_leaf_110_clk _00283_ VGND VGND VPWR VPWR _234_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12015_ _152_\[26\] _06007_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__or2_1
XFILLER_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13966_ clknet_leaf_97_clk _01185_ VGND VGND VPWR VPWR _118_\[14\] sky130_fd_sc_hd__dfxtp_2
X_13897_ clknet_leaf_64_clk _01116_ VGND VGND VPWR VPWR _122_\[9\] sky130_fd_sc_hd__dfxtp_1
X_12917_ clknet_leaf_88_clk _00141_ VGND VGND VPWR VPWR _116_\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12848_ _06468_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__clkbuf_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _06432_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09990_ _04157_ _04359_ _04360_ _04368_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__o31a_1
XFILLER_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08941_ _03296_ _03329_ _03330_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__or3_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08872_ _03290_ _03292_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07823_ _185_\[23\] _234_\[23\] VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__or2_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07754_ _182_\[21\] _01675_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__nand2_1
X_07685_ _02227_ _02229_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__xnor2_4
X_06705_ _118_\[17\] _116_\[17\] _01381_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__mux2_1
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06636_ _01304_ _01307_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_91_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_16
X_09424_ _03825_ _03826_ _03828_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__and3_1
XFILLER_52_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06567_ net35 _01253_ _01275_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__o21ai_4
X_09355_ _03722_ _03741_ _03761_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__o21ai_2
XFILLER_33_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06498_ net33 _01211_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__or2_2
X_08306_ _225_\[1\] VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__buf_4
X_09286_ _03693_ _03694_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__nand2_1
XFILLER_21_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08237_ _231_\[13\] _02690_ _02712_ _02722_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__a211o_1
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08168_ _167_\[26\] _02652_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__or2_1
XFILLER_69_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07119_ _240_\[25\] _01649_ _01607_ _01689_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__a211o_1
X_08099_ _01670_ _02623_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__or2_1
X_10130_ _01233_ _03978_ _04499_ _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__o31a_1
X_10061_ _04078_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__buf_2
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13820_ clknet_leaf_68_clk _01039_ VGND VGND VPWR VPWR _128_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13751_ clknet_leaf_67_clk _00970_ VGND VGND VPWR VPWR _132_\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_62_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10963_ _01424_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__buf_2
X_12702_ _06392_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13682_ clknet_leaf_77_clk _00901_ VGND VGND VPWR VPWR _136_\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10894_ _04682_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__buf_2
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12633_ _126_\[9\] _124_\[9\] _06346_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__mux2_1
XFILLER_71_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12564_ _128_\[8\] _126_\[8\] _06313_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__mux2_1
XFILLER_129_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11515_ _118_\[13\] _05556_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12495_ _130_\[7\] _128_\[7\] _06280_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__mux2_1
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11446_ _116_\[3\] _05494_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__and2_1
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11377_ _05433_ _05434_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__or2_1
X_10328_ _182_\[24\] _04654_ _04642_ _04650_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__a31o_1
X_13116_ clknet_leaf_119_clk _00335_ VGND VGND VPWR VPWR _231_\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13047_ clknet_leaf_109_clk _00266_ VGND VGND VPWR VPWR _237_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _01305_ _01338_ _04624_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__nor3_4
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13949_ clknet_leaf_90_clk _01168_ VGND VGND VPWR VPWR _120_\[29\] sky130_fd_sc_hd__dfxtp_1
X_07470_ _01989_ _01994_ _02021_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09140_ _02323_ _03524_ _03522_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__o21ai_1
X_09071_ _02262_ _03485_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__xnor2_1
X_08022_ _02516_ _02525_ _02554_ _01523_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__o31a_1
XFILLER_116_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09973_ _04351_ _04352_ _03945_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__a21o_1
XFILLER_104_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08924_ _02827_ _02787_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08855_ _03268_ _03269_ _03276_ _01439_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__o211a_1
X_07806_ _02341_ _02345_ _01354_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__o21a_1
X_08786_ _170_\[11\] _02804_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__and2_1
X_07737_ _02254_ _02279_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_64_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_53_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07668_ _02186_ _02206_ _02212_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__a21oi_1
XFILLER_41_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06619_ _392_\[1\] _01207_ _01209_ _01318_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__a31o_1
X_07599_ _02142_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__inv_2
XFILLER_71_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09407_ _02865_ _01884_ _03309_ _03812_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__a211o_1
X_09338_ _02868_ _03744_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11300_ _149_\[16\] _132_\[16\] VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__nand2_1
X_09269_ _02451_ _03677_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__xor2_1
X_12280_ _136_\[1\] _134_\[1\] _06167_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__mux2_1
XFILLER_119_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11231_ _05306_ _05307_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__nand2_1
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11162_ _05227_ _05249_ _05250_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__a21o_1
XFILLER_107_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10113_ _04484_ _04485_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__nor2_1
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11093_ _158_\[0\] _05193_ _05197_ _05198_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__a22o_1
XFILLER_122_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10044_ _01232_ _04415_ _04417_ _04420_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__a22o_1
XFILLER_76_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13803_ clknet_leaf_93_clk _01022_ VGND VGND VPWR VPWR _128_\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_55_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_16
X_11995_ _05909_ _05948_ _05988_ _05990_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__o31a_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13734_ clknet_leaf_59_clk _00953_ VGND VGND VPWR VPWR _132_\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10946_ net42 _05068_ _05104_ _05086_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__a211o_1
X_13665_ clknet_leaf_59_clk _00884_ VGND VGND VPWR VPWR _136_\[1\] sky130_fd_sc_hd__dfxtp_1
X_10877_ _167_\[27\] _05022_ _05043_ _05055_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__o211a_1
XFILLER_32_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12616_ _06347_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13596_ clknet_leaf_50_clk _00815_ VGND VGND VPWR VPWR _142_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12547_ _128_\[0\] _126_\[0\] _06302_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__mux2_1
XFILLER_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12478_ _132_\[31\] _130_\[31\] _06269_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__mux2_1
XANTENNA_3 _02293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11429_ _118_\[19\] _05479_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06970_ _01568_ _01576_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__or2_1
XFILLER_39_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08640_ _03065_ _03067_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_46_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_16
X_08571_ _02994_ _02999_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__nand2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07522_ _02071_ _02043_ _02042_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__o21a_1
XFILLER_34_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07453_ _01984_ _01985_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__or2b_1
XFILLER_50_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07384_ _01938_ _01939_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09123_ _03534_ _03535_ _03536_ _01523_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__o211a_1
XFILLER_135_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09054_ _03467_ _03468_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__or2b_1
X_08005_ _01629_ _01612_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__xnor2_2
XFILLER_116_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09956_ _01281_ _04087_ _04080_ _03938_ _04054_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__o311a_1
XFILLER_106_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09887_ _04266_ _04270_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__nand2_1
XFILLER_106_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ _228_\[15\] _231_\[15\] _03326_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__o21a_2
X_08838_ _02074_ _03259_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_37_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_73_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08769_ _185_\[11\] _03192_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11780_ _05792_ _05794_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__nand2_1
XFILLER_60_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10800_ _164_\[4\] _04986_ _05000_ _05001_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__a211o_1
XFILLER_53_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10731_ _167_\[16\] _04945_ _04951_ _04952_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__a211o_1
XFILLER_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13450_ clknet_leaf_3_clk _00669_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfxtp_2
XFILLER_13_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12401_ _132_\[26\] _134_\[26\] _06230_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__mux2_1
X_10662_ _173_\[28\] _04848_ _04903_ _04839_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__a211o_1
XFILLER_41_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10593_ _173_\[5\] _04849_ _04857_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__a21o_1
X_13381_ clknet_leaf_125_clk _00600_ VGND VGND VPWR VPWR _170_\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12332_ _136_\[26\] _134_\[26\] _06189_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__mux2_1
XFILLER_5_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12263_ _138_\[25\] _136_\[25\] _06156_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__mux2_1
XFILLER_5_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11214_ _149_\[5\] _132_\[5\] VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__or2_1
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12194_ _140_\[24\] _138_\[24\] _06123_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__mux2_1
XFILLER_107_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput51 net51 VGND VGND VPWR VPWR dout[23] sky130_fd_sc_hd__buf_2
Xoutput40 net40 VGND VGND VPWR VPWR dout[13] sky130_fd_sc_hd__buf_2
X_11145_ net15 _05202_ _05193_ _158_\[13\] VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__a22o_1
Xoutput62 net62 VGND VGND VPWR VPWR dout[4] sky130_fd_sc_hd__buf_2
X_11076_ _03841_ _04691_ _05187_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10027_ _04398_ _04404_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__and2_1
XFILLER_0_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_28_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_63_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11978_ _140_\[10\] _140_\[8\] VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__nand2_1
XFILLER_91_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13717_ clknet_leaf_77_clk _00936_ VGND VGND VPWR VPWR _134_\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10929_ _164_\[10\] _05059_ _05043_ _05092_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__o211a_1
XFILLER_31_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13648_ clknet_leaf_47_clk _00867_ VGND VGND VPWR VPWR _138_\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13579_ clknet_leaf_51_clk _00798_ VGND VGND VPWR VPWR _142_\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09810_ _04169_ _04170_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__and2b_1
XFILLER_87_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09741_ _246_\[9\] _01314_ _04129_ _243_\[9\] _01457_ VGND VGND VPWR VPWR _04130_
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06953_ _243_\[16\] _01536_ _01557_ _01564_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__a211o_1
XFILLER_100_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09672_ _142_\[5\] _04023_ _04035_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__a21bo_1
X_06884_ _01444_ _01514_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__nand2_1
XFILLER_82_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08623_ _02999_ _03020_ _03051_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08554_ _02949_ _02952_ _02984_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__o21ai_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07505_ _02054_ _02055_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__and2b_1
XFILLER_63_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08485_ _02915_ _02917_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__xor2_1
XFILLER_50_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07436_ _01986_ _01988_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__nand2_1
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07367_ _01408_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__clkbuf_8
XFILLER_136_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09106_ _02804_ _02776_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07298_ _01427_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__clkbuf_8
X_09037_ _03450_ _03452_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_13_0_clk clknet_3_6_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_09939_ _01243_ _03950_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__nand2_1
X_12950_ clknet_leaf_29_clk _00169_ VGND VGND VPWR VPWR _246_\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _06485_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__clkbuf_1
X_11901_ _152_\[16\] _05903_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__or2_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11832_ _05842_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11763_ _140_\[21\] _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__xnor2_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13502_ clknet_leaf_37_clk _00721_ VGND VGND VPWR VPWR _158_\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _05694_ _05717_ _05716_ _05699_ _05705_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__o221a_1
X_10714_ _173_\[12\] _04917_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__or2_1
XFILLER_14_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10645_ _02353_ _04892_ _04630_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__mux2_1
XFILLER_42_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13433_ clknet_leaf_123_clk _00652_ VGND VGND VPWR VPWR _164_\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13364_ clknet_leaf_124_clk _00583_ VGND VGND VPWR VPWR _170_\[14\] sky130_fd_sc_hd__dfxtp_1
X_12315_ _01393_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__clkbuf_4
X_10576_ _173_\[0\] _176_\[0\] _01226_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__mux2_1
XFILLER_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13295_ clknet_leaf_26_clk _00514_ VGND VGND VPWR VPWR _176_\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12246_ _138_\[17\] _136_\[17\] _06145_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__mux2_1
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12177_ _140_\[16\] _138_\[16\] _06112_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__mux2_1
XFILLER_69_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11128_ net10 _05190_ _05192_ _158_\[9\] VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__a22o_1
XFILLER_96_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11059_ _164_\[24\] _01218_ _04648_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__o21a_1
XFILLER_37_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08270_ _02686_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__or2_1
X_07221_ _185_\[3\] _234_\[3\] VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__nand2_1
XFILLER_32_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07152_ _185_\[0\] _234_\[0\] VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__or2_1
XFILLER_145_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07083_ _173_\[17\] _01661_ _01617_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_8_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_133_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07985_ _02468_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__inv_2
X_09724_ _142_\[8\] _04113_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__and2_1
X_06936_ _243_\[11\] _01536_ _01509_ _01552_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__a211o_1
XFILLER_55_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09655_ _142_\[6\] _04045_ _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__and3_1
X_06867_ _246_\[24\] _01496_ _01460_ _01502_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__a211o_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08606_ _02862_ _03034_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__xnor2_2
X_09586_ _01241_ _03925_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__nand2_1
X_06798_ _246_\[6\] _01422_ _01425_ _01451_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__o211a_1
Xclkbuf_3_2_0_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _02967_ _02964_ _02965_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__nor3_1
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08468_ _228_\[1\] _231_\[1\] _02901_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__o21a_1
X_07419_ _01632_ _01827_ _01693_ _01972_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__a211o_1
XFILLER_109_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10430_ _176_\[21\] _04735_ _04742_ _04740_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__o211a_1
X_08399_ _02842_ _01801_ _02824_ _02843_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__o211a_1
XFILLER_136_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10361_ _01214_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__buf_4
X_12100_ _06076_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__clkbuf_1
X_10292_ _01417_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13080_ clknet_leaf_100_clk _00299_ VGND VGND VPWR VPWR _234_\[24\] sky130_fd_sc_hd__dfxtp_1
X_12031_ _06022_ _06023_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13982_ clknet_leaf_68_clk _01201_ VGND VGND VPWR VPWR _118_\[30\] sky130_fd_sc_hd__dfxtp_2
XFILLER_93_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12933_ clknet_leaf_39_clk _00152_ VGND VGND VPWR VPWR _246_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _118_\[23\] _120_\[23\] _06473_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__mux2_1
XFILLER_18_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _05793_ _05806_ _05801_ _05826_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__o31a_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12795_ _122_\[22\] _120_\[22\] _06434_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__mux2_1
X_11746_ net23 _05763_ _05742_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__mux2_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11677_ _05702_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10628_ _176_\[17\] _04684_ _01417_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__a21o_1
X_13416_ clknet_leaf_1_clk _00635_ VGND VGND VPWR VPWR _164_\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10559_ _179_\[27\] _04799_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__or2_1
XFILLER_6_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13347_ clknet_leaf_4_clk _00566_ VGND VGND VPWR VPWR _173_\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13278_ clknet_leaf_7_clk _00497_ VGND VGND VPWR VPWR _179_\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12229_ _138_\[9\] _136_\[9\] _06134_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__mux2_1
XFILLER_130_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07770_ _02310_ _02311_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__xnor2_1
X_06721_ _01393_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__buf_4
XFILLER_65_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09440_ _03762_ _03765_ _03800_ _03802_ _03834_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__a311o_1
XFILLER_25_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06652_ _01295_ _01252_ _01326_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__a21o_1
XFILLER_64_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06583_ _01276_ _01285_ _01244_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__a21oi_1
X_09371_ _03758_ _03760_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__and2b_1
X_08322_ _225_\[5\] VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__clkbuf_4
X_08253_ _164_\[18\] _02701_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__or2_1
XFILLER_138_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07204_ _01736_ _01764_ _01765_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__and3_1
XFILLER_118_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08184_ _167_\[31\] _02652_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__or2_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07135_ _173_\[29\] _01701_ _01672_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__mux2_1
XFILLER_134_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07066_ _240_\[13\] _01583_ _01607_ _01648_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__a211o_1
XFILLER_145_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07968_ _01694_ _02448_ _02419_ _02503_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__o211a_1
X_09707_ _04095_ _04097_ _03867_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__o21ai_1
X_06919_ _243_\[6\] _01485_ _01481_ _01540_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__o211a_1
XFILLER_75_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07899_ _02396_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__inv_2
XFILLER_28_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09638_ _01280_ _03896_ _03950_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__o21ai_1
XFILLER_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09569_ _246_\[2\] _01313_ _03913_ _243_\[2\] _01432_ VGND VGND VPWR VPWR _03965_
+ sky130_fd_sc_hd__o221a_1
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11600_ _05631_ _05633_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__or2_1
X_12580_ _06328_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11531_ _05570_ _05571_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11462_ _118_\[23\] _118_\[12\] VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__xnor2_1
X_13201_ clknet_leaf_35_clk _00420_ VGND VGND VPWR VPWR _185_\[11\] sky130_fd_sc_hd__dfxtp_2
X_11393_ _05409_ _05414_ _05422_ _05448_ _05416_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__o311a_1
X_10413_ _176_\[16\] _04725_ _04730_ _04728_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__a211o_1
X_10344_ _179_\[30\] _04658_ _04679_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__a21o_1
X_13132_ clknet_leaf_109_clk _00351_ VGND VGND VPWR VPWR _228_\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10275_ _182_\[1\] _04634_ _04639_ _00105_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__o211a_1
X_13063_ clknet_leaf_109_clk _00282_ VGND VGND VPWR VPWR _234_\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ _152_\[26\] _06007_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__nand2_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13965_ clknet_leaf_97_clk _01184_ VGND VGND VPWR VPWR _118_\[13\] sky130_fd_sc_hd__dfxtp_2
X_13896_ clknet_leaf_64_clk _01115_ VGND VGND VPWR VPWR _122_\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12916_ clknet_leaf_88_clk _00140_ VGND VGND VPWR VPWR _116_\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12847_ _118_\[15\] _120_\[15\] _06462_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__mux2_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _122_\[14\] _120_\[14\] _06423_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__mux2_1
X_11729_ _142_\[0\] _05748_ _05625_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__mux2_1
XFILLER_128_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08940_ _03357_ _03358_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__xnor2_2
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08871_ _228_\[14\] _231_\[14\] _03291_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__o21a_1
XFILLER_84_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07822_ _01701_ _02361_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__xnor2_2
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07753_ _01671_ _01973_ _01886_ _02295_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__o211a_1
X_07684_ _182_\[17\] _01661_ _02173_ _02228_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__o22a_2
X_06704_ _01384_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06635_ _01298_ _01305_ _01320_ _01337_ VGND VGND VPWR VPWR _436_\[0\] sky130_fd_sc_hd__a211o_1
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09423_ _228_\[30\] _231_\[30\] _03827_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__o21a_1
XFILLER_25_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09354_ _03758_ _03760_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__xnor2_1
X_06566_ net35 _01271_ _01272_ _01274_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__o211a_1
XFILLER_52_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08305_ _01799_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__clkbuf_4
X_06497_ _01206_ _01210_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__or2_1
X_09285_ _03660_ _03657_ _03658_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__a21bo_1
XFILLER_60_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08236_ _228_\[13\] _02698_ _02679_ _02721_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__o211a_1
X_08167_ _234_\[25\] _02659_ _02636_ _02672_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__o211a_1
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07118_ _01687_ _01639_ _01609_ _01688_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__o211a_1
XFILLER_4_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08098_ _167_\[6\] _231_\[6\] _01672_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__mux2_1
XFILLER_133_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07049_ _237_\[10\] VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__buf_4
XFILLER_133_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10060_ _01284_ _04005_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__nand2_1
XFILLER_88_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13750_ clknet_leaf_67_clk _00969_ VGND VGND VPWR VPWR _132_\[22\] sky130_fd_sc_hd__dfxtp_2
XFILLER_90_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10962_ _05079_ _05115_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__or2_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12701_ _124_\[9\] _122_\[9\] _06390_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__mux2_1
XFILLER_83_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13681_ clknet_leaf_78_clk _00900_ VGND VGND VPWR VPWR _136_\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10893_ _164_\[31\] _05048_ _05066_ _05067_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__o211a_1
XFILLER_16_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12632_ _06355_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12563_ _06319_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12494_ _06283_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11514_ _118_\[28\] _118_\[17\] VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11445_ _118_\[21\] _05493_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11376_ _149_\[26\] _132_\[26\] VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__and2_1
XFILLER_125_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10327_ _179_\[23\] _04658_ _04669_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__a21o_1
X_13115_ clknet_leaf_120_clk _00334_ VGND VGND VPWR VPWR _231_\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _01272_ _01349_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__nand2_1
XFILLER_105_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13046_ clknet_leaf_108_clk _00265_ VGND VGND VPWR VPWR _237_\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10189_ _142_\[28\] _04557_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__nor2_1
XFILLER_94_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13948_ clknet_leaf_89_clk _01167_ VGND VGND VPWR VPWR _120_\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13879_ clknet_leaf_92_clk _01098_ VGND VGND VPWR VPWR _124_\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09070_ _185_\[20\] _03484_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__xor2_1
X_08021_ _02516_ _02525_ _02554_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__o21ai_1
XFILLER_128_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09972_ _04347_ _04350_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__or2_1
XFILLER_104_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08923_ _02117_ _03315_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__or2_1
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08854_ _02404_ _03275_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__nand2_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08785_ _03187_ _03188_ _03207_ _01923_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__a31o_1
X_07805_ _02341_ _02345_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__nand2_1
X_07736_ _02218_ _02255_ _02276_ _02222_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__o22ai_1
XFILLER_38_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07667_ _02208_ _02211_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__xor2_1
X_06618_ _01251_ _01209_ _01273_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__and3b_1
X_07598_ _02052_ _02078_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__nand2_1
XFILLER_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09406_ _01409_ _03804_ _03805_ _03811_ _01799_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__o311a_1
XFILLER_25_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06549_ _158_\[9\] _01257_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__or2_1
XFILLER_40_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09337_ _02827_ _02797_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09268_ _185_\[26\] _03676_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__xnor2_1
X_08219_ _228_\[8\] _02698_ _02679_ _02709_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__o211a_1
XFILLER_119_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09199_ _02362_ _03609_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__nand2_1
X_11230_ _149_\[7\] _132_\[7\] VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__nand2_1
XFILLER_106_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11161_ net19 _05202_ _05193_ _158_\[17\] VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__a22o_1
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10112_ _04484_ _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__and2_1
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11092_ net32 _05196_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__or2_1
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10043_ _01232_ _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__nor2_1
XFILLER_75_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13802_ clknet_leaf_86_clk _01021_ VGND VGND VPWR VPWR _128_\[10\] sky130_fd_sc_hd__dfxtp_1
X_11994_ _05966_ _05976_ _05977_ _05989_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__o211a_1
XFILLER_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13733_ clknet_leaf_61_clk _00952_ VGND VGND VPWR VPWR _132_\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10945_ _164_\[15\] _05059_ _05094_ _05103_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__o211a_1
X_13664_ clknet_leaf_58_clk _00883_ VGND VGND VPWR VPWR _136_\[0\] sky130_fd_sc_hd__dfxtp_1
X_10876_ _170_\[27\] _05036_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__or2_1
X_12615_ _126_\[0\] _124_\[0\] _06346_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__mux2_1
XFILLER_129_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13595_ clknet_leaf_50_clk _00814_ VGND VGND VPWR VPWR _142_\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12546_ _06310_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12477_ _06274_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11428_ _118_\[8\] _118_\[4\] VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__xnor2_1
XANTENNA_4 _02353_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11359_ _05263_ _05419_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__nand2_1
XFILLER_99_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13029_ clknet_leaf_42_clk _00248_ VGND VGND VPWR VPWR _237_\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08570_ _02781_ _02845_ _02834_ _03000_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__o211a_1
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07521_ _02040_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__inv_2
XFILLER_47_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07452_ _01635_ _01973_ _01886_ _02004_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__o211a_1
XFILLER_23_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07383_ _243_\[8\] _240_\[8\] _01629_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__mux2_4
XFILLER_50_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09122_ _03534_ _03535_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__nand2_1
X_09053_ _170_\[20\] _02835_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__nand2_1
XFILLER_144_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08004_ _02513_ _02514_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__and2b_1
XFILLER_143_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09955_ _01237_ _03876_ _04083_ _04334_ _01231_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__o311a_1
XFILLER_89_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09886_ _04205_ _04267_ _04269_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__o21a_1
XFILLER_106_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08906_ _228_\[15\] _231_\[15\] _02817_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__a21o_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08837_ _03256_ _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__xor2_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08768_ _02849_ _03191_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__xnor2_2
XFILLER_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07719_ _01707_ _02261_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__xnor2_4
X_08699_ _01778_ _03125_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__nor2_1
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10730_ _01418_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__clkbuf_4
X_10661_ _176_\[28\] _04872_ _04633_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__o211a_1
X_12400_ _06234_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__clkbuf_1
X_10592_ _176_\[5\] net68 _01833_ _04692_ _02711_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__a221o_1
X_13380_ clknet_leaf_128_clk _00599_ VGND VGND VPWR VPWR _170_\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12331_ _06197_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12262_ _06161_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11213_ _05292_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12193_ _06125_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__clkbuf_1
Xoutput41 net41 VGND VGND VPWR VPWR dout[14] sky130_fd_sc_hd__buf_2
Xoutput52 net52 VGND VGND VPWR VPWR dout[24] sky130_fd_sc_hd__buf_2
X_11144_ _158_\[13\] _01260_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__xnor2_1
Xoutput63 net63 VGND VGND VPWR VPWR dout[5] sky130_fd_sc_hd__buf_2
XFILLER_1_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11075_ _164_\[30\] _01226_ _04637_ net59 _01417_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__a221o_1
XFILLER_1_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10026_ _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__inv_2
XFILLER_76_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11977_ _140_\[10\] _140_\[8\] VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__or2_1
XFILLER_91_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13716_ clknet_leaf_77_clk _00935_ VGND VGND VPWR VPWR _134_\[20\] sky130_fd_sc_hd__dfxtp_1
X_10928_ _167_\[10\] _05089_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__or2_1
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13647_ clknet_leaf_47_clk _00866_ VGND VGND VPWR VPWR _138_\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10859_ _04685_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__buf_2
X_13578_ clknet_leaf_35_clk _00797_ VGND VGND VPWR VPWR _142_\[10\] sky130_fd_sc_hd__dfxtp_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12529_ _06301_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09740_ _03914_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__buf_2
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06952_ _240_\[16\] _01526_ _01558_ _01563_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__o211a_1
.ends

