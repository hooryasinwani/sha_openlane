magic
tech sky130A
magscale 1 2
timestamp 1733415340
<< obsli1 >>
rect 1104 2159 80592 81617
<< obsm1 >>
rect 14 1640 81222 81648
<< metal2 >>
rect 3238 83088 3294 83688
rect 7746 83088 7802 83688
rect 12254 83088 12310 83688
rect 16762 83088 16818 83688
rect 21270 83088 21326 83688
rect 25778 83088 25834 83688
rect 30930 83088 30986 83688
rect 35438 83088 35494 83688
rect 39946 83088 40002 83688
rect 44454 83088 44510 83688
rect 48962 83088 49018 83688
rect 53470 83088 53526 83688
rect 58622 83088 58678 83688
rect 63130 83088 63186 83688
rect 67638 83088 67694 83688
rect 72146 83088 72202 83688
rect 76654 83088 76710 83688
rect 81162 83088 81218 83688
rect 18 200 74 800
rect 4526 200 4582 800
rect 9034 200 9090 800
rect 13542 200 13598 800
rect 18050 200 18106 800
rect 22558 200 22614 800
rect 27710 200 27766 800
rect 32218 200 32274 800
rect 36726 200 36782 800
rect 41234 200 41290 800
rect 45742 200 45798 800
rect 50250 200 50306 800
rect 55402 200 55458 800
rect 59910 200 59966 800
rect 64418 200 64474 800
rect 68926 200 68982 800
rect 73434 200 73490 800
rect 77942 200 77998 800
<< obsm2 >>
rect 20 83032 3182 83178
rect 3350 83032 7690 83178
rect 7858 83032 12198 83178
rect 12366 83032 16706 83178
rect 16874 83032 21214 83178
rect 21382 83032 25722 83178
rect 25890 83032 30874 83178
rect 31042 83032 35382 83178
rect 35550 83032 39890 83178
rect 40058 83032 44398 83178
rect 44566 83032 48906 83178
rect 49074 83032 53414 83178
rect 53582 83032 58566 83178
rect 58734 83032 63074 83178
rect 63242 83032 67582 83178
rect 67750 83032 72090 83178
rect 72258 83032 76598 83178
rect 76766 83032 81106 83178
rect 20 856 81216 83032
rect 130 734 4470 856
rect 4638 734 8978 856
rect 9146 734 13486 856
rect 13654 734 17994 856
rect 18162 734 22502 856
rect 22670 734 27654 856
rect 27822 734 32162 856
rect 32330 734 36670 856
rect 36838 734 41178 856
rect 41346 734 45686 856
rect 45854 734 50194 856
rect 50362 734 55346 856
rect 55514 734 59854 856
rect 60022 734 64362 856
rect 64530 734 68870 856
rect 69038 734 73378 856
rect 73546 734 77886 856
rect 78054 734 81216 856
<< metal3 >>
rect 200 82288 800 82408
rect 80944 78888 81544 79008
rect 200 77528 800 77648
rect 80944 74128 81544 74248
rect 200 72768 800 72888
rect 80944 69368 81544 69488
rect 200 68008 800 68128
rect 80944 64608 81544 64728
rect 200 63248 800 63368
rect 80944 59848 81544 59968
rect 200 58488 800 58608
rect 80944 54408 81544 54528
rect 200 53048 800 53168
rect 80944 49648 81544 49768
rect 200 48288 800 48408
rect 80944 44888 81544 45008
rect 200 43528 800 43648
rect 80944 40128 81544 40248
rect 200 38768 800 38888
rect 80944 35368 81544 35488
rect 200 34008 800 34128
rect 80944 30608 81544 30728
rect 200 29248 800 29368
rect 80944 25168 81544 25288
rect 200 23808 800 23928
rect 80944 20408 81544 20528
rect 200 19048 800 19168
rect 80944 15648 81544 15768
rect 200 14288 800 14408
rect 80944 10888 81544 11008
rect 200 9528 800 9648
rect 80944 6128 81544 6248
rect 200 4768 800 4888
rect 80944 1368 81544 1488
<< obsm3 >>
rect 880 82208 80944 82381
rect 800 79088 80944 82208
rect 800 78808 80864 79088
rect 800 77728 80944 78808
rect 880 77448 80944 77728
rect 800 74328 80944 77448
rect 800 74048 80864 74328
rect 800 72968 80944 74048
rect 880 72688 80944 72968
rect 800 69568 80944 72688
rect 800 69288 80864 69568
rect 800 68208 80944 69288
rect 880 67928 80944 68208
rect 800 64808 80944 67928
rect 800 64528 80864 64808
rect 800 63448 80944 64528
rect 880 63168 80944 63448
rect 800 60048 80944 63168
rect 800 59768 80864 60048
rect 800 58688 80944 59768
rect 880 58408 80944 58688
rect 800 54608 80944 58408
rect 800 54328 80864 54608
rect 800 53248 80944 54328
rect 880 52968 80944 53248
rect 800 49848 80944 52968
rect 800 49568 80864 49848
rect 800 48488 80944 49568
rect 880 48208 80944 48488
rect 800 45088 80944 48208
rect 800 44808 80864 45088
rect 800 43728 80944 44808
rect 880 43448 80944 43728
rect 800 40328 80944 43448
rect 800 40048 80864 40328
rect 800 38968 80944 40048
rect 880 38688 80944 38968
rect 800 35568 80944 38688
rect 800 35288 80864 35568
rect 800 34208 80944 35288
rect 880 33928 80944 34208
rect 800 30808 80944 33928
rect 800 30528 80864 30808
rect 800 29448 80944 30528
rect 880 29168 80944 29448
rect 800 25368 80944 29168
rect 800 25088 80864 25368
rect 800 24008 80944 25088
rect 880 23728 80944 24008
rect 800 20608 80944 23728
rect 800 20328 80864 20608
rect 800 19248 80944 20328
rect 880 18968 80944 19248
rect 800 15848 80944 18968
rect 800 15568 80864 15848
rect 800 14488 80944 15568
rect 880 14208 80944 14488
rect 800 11088 80944 14208
rect 800 10808 80864 11088
rect 800 9728 80944 10808
rect 880 9448 80944 9728
rect 800 6328 80944 9448
rect 800 6048 80864 6328
rect 800 4968 80944 6048
rect 880 4688 80944 4968
rect 800 1568 80944 4688
rect 800 1395 80864 1568
<< metal4 >>
rect 4208 2128 4528 81648
rect 4868 2128 5188 81648
rect 34928 2128 35248 81648
rect 35588 2128 35908 81648
rect 65648 2128 65968 81648
rect 66308 2128 66628 81648
<< obsm4 >>
rect 1899 2211 4128 81293
rect 4608 2211 4788 81293
rect 5268 2211 34848 81293
rect 35328 2211 35508 81293
rect 35988 2211 65568 81293
rect 66048 2211 66228 81293
rect 66708 2211 79981 81293
<< metal5 >>
rect 1056 67278 80640 67598
rect 1056 66618 80640 66938
rect 1056 36642 80640 36962
rect 1056 35982 80640 36302
rect 1056 6006 80640 6326
rect 1056 5346 80640 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 81648 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 81648 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 81648 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 80640 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 80640 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67278 80640 67598 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 81648 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 81648 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 81648 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 80640 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 80640 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 80640 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 18050 200 18106 800 6 clk
port 3 nsew signal input
rlabel metal3 s 80944 35368 81544 35488 6 din[0]
port 4 nsew signal input
rlabel metal3 s 200 72768 800 72888 6 din[10]
port 5 nsew signal input
rlabel metal2 s 59910 200 59966 800 6 din[11]
port 6 nsew signal input
rlabel metal2 s 7746 83088 7802 83688 6 din[12]
port 7 nsew signal input
rlabel metal3 s 80944 54408 81544 54528 6 din[13]
port 8 nsew signal input
rlabel metal2 s 77942 200 77998 800 6 din[14]
port 9 nsew signal input
rlabel metal3 s 80944 10888 81544 11008 6 din[15]
port 10 nsew signal input
rlabel metal3 s 80944 15648 81544 15768 6 din[16]
port 11 nsew signal input
rlabel metal3 s 200 19048 800 19168 6 din[17]
port 12 nsew signal input
rlabel metal3 s 80944 64608 81544 64728 6 din[18]
port 13 nsew signal input
rlabel metal3 s 200 82288 800 82408 6 din[19]
port 14 nsew signal input
rlabel metal3 s 80944 59848 81544 59968 6 din[1]
port 15 nsew signal input
rlabel metal3 s 80944 6128 81544 6248 6 din[20]
port 16 nsew signal input
rlabel metal2 s 25778 83088 25834 83688 6 din[21]
port 17 nsew signal input
rlabel metal3 s 80944 25168 81544 25288 6 din[22]
port 18 nsew signal input
rlabel metal2 s 27710 200 27766 800 6 din[23]
port 19 nsew signal input
rlabel metal3 s 200 48288 800 48408 6 din[24]
port 20 nsew signal input
rlabel metal3 s 80944 49648 81544 49768 6 din[25]
port 21 nsew signal input
rlabel metal2 s 68926 200 68982 800 6 din[26]
port 22 nsew signal input
rlabel metal3 s 200 68008 800 68128 6 din[27]
port 23 nsew signal input
rlabel metal2 s 45742 200 45798 800 6 din[28]
port 24 nsew signal input
rlabel metal3 s 200 58488 800 58608 6 din[29]
port 25 nsew signal input
rlabel metal2 s 36726 200 36782 800 6 din[2]
port 26 nsew signal input
rlabel metal2 s 35438 83088 35494 83688 6 din[30]
port 27 nsew signal input
rlabel metal2 s 63130 83088 63186 83688 6 din[31]
port 28 nsew signal input
rlabel metal2 s 16762 83088 16818 83688 6 din[3]
port 29 nsew signal input
rlabel metal3 s 200 63248 800 63368 6 din[4]
port 30 nsew signal input
rlabel metal3 s 200 38768 800 38888 6 din[5]
port 31 nsew signal input
rlabel metal2 s 81162 83088 81218 83688 6 din[6]
port 32 nsew signal input
rlabel metal2 s 73434 200 73490 800 6 din[7]
port 33 nsew signal input
rlabel metal2 s 44454 83088 44510 83688 6 din[8]
port 34 nsew signal input
rlabel metal3 s 80944 78888 81544 79008 6 din[9]
port 35 nsew signal input
rlabel metal2 s 64418 200 64474 800 6 dout[0]
port 36 nsew signal output
rlabel metal2 s 39946 83088 40002 83688 6 dout[10]
port 37 nsew signal output
rlabel metal3 s 200 9528 800 9648 6 dout[11]
port 38 nsew signal output
rlabel metal3 s 80944 20408 81544 20528 6 dout[12]
port 39 nsew signal output
rlabel metal2 s 50250 200 50306 800 6 dout[13]
port 40 nsew signal output
rlabel metal3 s 80944 30608 81544 30728 6 dout[14]
port 41 nsew signal output
rlabel metal2 s 53470 83088 53526 83688 6 dout[15]
port 42 nsew signal output
rlabel metal2 s 58622 83088 58678 83688 6 dout[16]
port 43 nsew signal output
rlabel metal2 s 3238 83088 3294 83688 6 dout[17]
port 44 nsew signal output
rlabel metal2 s 18 200 74 800 6 dout[18]
port 45 nsew signal output
rlabel metal3 s 200 53048 800 53168 6 dout[19]
port 46 nsew signal output
rlabel metal2 s 48962 83088 49018 83688 6 dout[1]
port 47 nsew signal output
rlabel metal3 s 200 34008 800 34128 6 dout[20]
port 48 nsew signal output
rlabel metal3 s 200 14288 800 14408 6 dout[21]
port 49 nsew signal output
rlabel metal2 s 30930 83088 30986 83688 6 dout[22]
port 50 nsew signal output
rlabel metal2 s 9034 200 9090 800 6 dout[23]
port 51 nsew signal output
rlabel metal2 s 4526 200 4582 800 6 dout[24]
port 52 nsew signal output
rlabel metal3 s 80944 74128 81544 74248 6 dout[25]
port 53 nsew signal output
rlabel metal2 s 76654 83088 76710 83688 6 dout[26]
port 54 nsew signal output
rlabel metal2 s 32218 200 32274 800 6 dout[27]
port 55 nsew signal output
rlabel metal3 s 80944 69368 81544 69488 6 dout[28]
port 56 nsew signal output
rlabel metal3 s 80944 1368 81544 1488 6 dout[29]
port 57 nsew signal output
rlabel metal3 s 200 23808 800 23928 6 dout[2]
port 58 nsew signal output
rlabel metal3 s 200 4768 800 4888 6 dout[30]
port 59 nsew signal output
rlabel metal2 s 13542 200 13598 800 6 dout[31]
port 60 nsew signal output
rlabel metal2 s 22558 200 22614 800 6 dout[3]
port 61 nsew signal output
rlabel metal3 s 200 43528 800 43648 6 dout[4]
port 62 nsew signal output
rlabel metal3 s 80944 44888 81544 45008 6 dout[5]
port 63 nsew signal output
rlabel metal2 s 41234 200 41290 800 6 dout[6]
port 64 nsew signal output
rlabel metal2 s 72146 83088 72202 83688 6 dout[7]
port 65 nsew signal output
rlabel metal2 s 67638 83088 67694 83688 6 dout[8]
port 66 nsew signal output
rlabel metal2 s 12254 83088 12310 83688 6 dout[9]
port 67 nsew signal output
rlabel metal2 s 21270 83088 21326 83688 6 dst_ready
port 68 nsew signal input
rlabel metal2 s 55402 200 55458 800 6 dst_write
port 69 nsew signal output
rlabel metal3 s 200 29248 800 29368 6 rst
port 70 nsew signal input
rlabel metal3 s 200 77528 800 77648 6 src_read
port 71 nsew signal output
rlabel metal3 s 80944 40128 81544 40248 6 src_ready
port 72 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 81744 83888
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 22013518
string GDS_FILE /openlane/designs/sha256/runs/RUN_2024.12.05_16.00.43/results/signoff/sha2_top.magic.gds
string GDS_START 1014022
<< end >>

